vram[12'h000] = 8'h1c;
vram[12'h001] = 8'h1d;
vram[12'h002] = 8'h1c;
vram[12'h003] = 8'h1d;
vram[12'h004] = 8'h1c;
vram[12'h005] = 8'h1d;
vram[12'h006] = 8'h1c;
vram[12'h007] = 8'h1d;
vram[12'h008] = 8'h1c;
vram[12'h009] = 8'h1d;
vram[12'h00a] = 8'h1c;
vram[12'h00b] = 8'h1d;
vram[12'h00c] = 8'h1c;
vram[12'h00d] = 8'h1d;
vram[12'h00e] = 8'h1c;
vram[12'h00f] = 8'h1d;
vram[12'h010] = 8'h1c;
vram[12'h011] = 8'h1d;
vram[12'h012] = 8'h1c;
vram[12'h013] = 8'h1d;
vram[12'h014] = 8'h1c;
vram[12'h015] = 8'h1d;
vram[12'h016] = 8'h1c;
vram[12'h017] = 8'h1d;
vram[12'h018] = 8'h1c;
vram[12'h019] = 8'h1d;
vram[12'h01a] = 8'h1c;
vram[12'h01b] = 8'h1d;
vram[12'h01c] = 8'h1c;
vram[12'h01d] = 8'h1d;
vram[12'h01e] = 8'h1c;
vram[12'h01f] = 8'h1d;
vram[12'h020] = 8'h20;
vram[12'h021] = 8'h20;
vram[12'h022] = 8'h20;
vram[12'h023] = 8'h20;
vram[12'h024] = 8'h20;
vram[12'h025] = 8'h20;
vram[12'h026] = 8'h20;
vram[12'h027] = 8'h20;
vram[12'h028] = 8'h20;
vram[12'h029] = 8'h20;
vram[12'h02a] = 8'h20;
vram[12'h02b] = 8'h20;
vram[12'h02c] = 8'h20;
vram[12'h02d] = 8'h20;
vram[12'h02e] = 8'h20;
vram[12'h02f] = 8'h20;
vram[12'h030] = 8'h20;
vram[12'h031] = 8'h20;
vram[12'h032] = 8'h20;
vram[12'h033] = 8'h20;
vram[12'h034] = 8'h20;
vram[12'h035] = 8'h20;
vram[12'h036] = 8'h20;
vram[12'h037] = 8'h20;
vram[12'h038] = 8'h20;
vram[12'h039] = 8'h20;
vram[12'h03a] = 8'h20;
vram[12'h03b] = 8'h20;
vram[12'h03c] = 8'h20;
vram[12'h03d] = 8'h20;
vram[12'h03e] = 8'h20;
vram[12'h03f] = 8'h54;
vram[12'h040] = 8'h69;
vram[12'h041] = 8'h6e;
vram[12'h042] = 8'h79;
vram[12'h043] = 8'h36;
vram[12'h044] = 8'h35;
vram[12'h045] = 8'h30;
vram[12'h046] = 8'h32;
vram[12'h047] = 8'h20;
vram[12'h048] = 8'h61;
vram[12'h049] = 8'h6e;
vram[12'h04a] = 8'h64;
vram[12'h04b] = 8'h20;
vram[12'h04c] = 8'h54;
vram[12'h04d] = 8'h69;
vram[12'h04e] = 8'h6e;
vram[12'h04f] = 8'h79;
vram[12'h050] = 8'h56;
vram[12'h051] = 8'h47;
vram[12'h052] = 8'h41;
vram[12'h053] = 8'h20;
vram[12'h054] = 8'h44;
vram[12'h055] = 8'h69;
vram[12'h056] = 8'h73;
vram[12'h057] = 8'h70;
vram[12'h058] = 8'h6c;
vram[12'h059] = 8'h61;
vram[12'h05a] = 8'h79;
vram[12'h05b] = 8'h20;
vram[12'h05c] = 8'h20;
vram[12'h05d] = 8'h20;
vram[12'h05e] = 8'h62;
vram[12'h05f] = 8'h79;
vram[12'h060] = 8'h20;
vram[12'h061] = 8'h43;
vram[12'h062] = 8'h46;
vram[12'h063] = 8'h32;
vram[12'h064] = 8'h30;
vram[12'h065] = 8'h37;
vram[12'h066] = 8'h2e;
vram[12'h067] = 8'h20;
vram[12'h068] = 8'h20;
vram[12'h069] = 8'h20;
vram[12'h06a] = 8'h20;
vram[12'h06b] = 8'h20;
vram[12'h06c] = 8'h20;
vram[12'h06d] = 8'h20;
vram[12'h06e] = 8'h20;
vram[12'h06f] = 8'h20;
vram[12'h070] = 8'h20;
vram[12'h071] = 8'h20;
vram[12'h072] = 8'h20;
vram[12'h073] = 8'h20;
vram[12'h074] = 8'h20;
vram[12'h075] = 8'h20;
vram[12'h076] = 8'h20;
vram[12'h077] = 8'h20;
vram[12'h078] = 8'h20;
vram[12'h079] = 8'h20;
vram[12'h07a] = 8'h20;
vram[12'h07b] = 8'h20;
vram[12'h07c] = 8'h20;
vram[12'h07d] = 8'h00;
vram[12'h07e] = 8'h00;
vram[12'h07f] = 8'h00;
vram[12'h080] = 8'h00;
vram[12'h081] = 8'h00;
vram[12'h082] = 8'h00;
vram[12'h083] = 8'h00;
vram[12'h084] = 8'h00;
vram[12'h085] = 8'h00;
vram[12'h086] = 8'h00;
vram[12'h087] = 8'h00;
vram[12'h088] = 8'h00;
vram[12'h089] = 8'h00;
vram[12'h08a] = 8'h00;
vram[12'h08b] = 8'h00;
vram[12'h08c] = 8'h00;
vram[12'h08d] = 8'h00;
vram[12'h08e] = 8'h00;
vram[12'h08f] = 8'h00;
vram[12'h090] = 8'h00;
vram[12'h091] = 8'h00;
vram[12'h092] = 8'h00;
vram[12'h093] = 8'h00;
vram[12'h094] = 8'h00;
vram[12'h095] = 8'h00;
vram[12'h096] = 8'h00;
vram[12'h097] = 8'h00;
vram[12'h098] = 8'h00;
vram[12'h099] = 8'h00;
vram[12'h09a] = 8'h00;
vram[12'h09b] = 8'h00;
vram[12'h09c] = 8'h00;
vram[12'h09d] = 8'h00;
vram[12'h09e] = 8'h00;
vram[12'h09f] = 8'h00;
vram[12'h0a0] = 8'h00;
vram[12'h0a1] = 8'h00;
vram[12'h0a2] = 8'h00;
vram[12'h0a3] = 8'h00;
vram[12'h0a4] = 8'h00;
vram[12'h0a5] = 8'h00;
vram[12'h0a6] = 8'h00;
vram[12'h0a7] = 8'h00;
vram[12'h0a8] = 8'h00;
vram[12'h0a9] = 8'h00;
vram[12'h0aa] = 8'h00;
vram[12'h0ab] = 8'h00;
vram[12'h0ac] = 8'h00;
vram[12'h0ad] = 8'h00;
vram[12'h0ae] = 8'h00;
vram[12'h0af] = 8'h00;
vram[12'h0b0] = 8'h00;
vram[12'h0b1] = 8'h00;
vram[12'h0b2] = 8'h00;
vram[12'h0b3] = 8'h00;
vram[12'h0b4] = 8'h00;
vram[12'h0b5] = 8'h00;
vram[12'h0b6] = 8'h00;
vram[12'h0b7] = 8'h00;
vram[12'h0b8] = 8'h00;
vram[12'h0b9] = 8'h00;
vram[12'h0ba] = 8'h00;
vram[12'h0bb] = 8'h00;
vram[12'h0bc] = 8'h00;
vram[12'h0bd] = 8'h00;
vram[12'h0be] = 8'h00;
vram[12'h0bf] = 8'h00;
vram[12'h0c0] = 8'h00;
vram[12'h0c1] = 8'h00;
vram[12'h0c2] = 8'h00;
vram[12'h0c3] = 8'h00;
vram[12'h0c4] = 8'h00;
vram[12'h0c5] = 8'h00;
vram[12'h0c6] = 8'h00;
vram[12'h0c7] = 8'h00;
vram[12'h0c8] = 8'h00;
vram[12'h0c9] = 8'h00;
vram[12'h0ca] = 8'h00;
vram[12'h0cb] = 8'h00;
vram[12'h0cc] = 8'h00;
vram[12'h0cd] = 8'h00;
vram[12'h0ce] = 8'h00;
vram[12'h0cf] = 8'h00;
vram[12'h0d0] = 8'h00;
vram[12'h0d1] = 8'h00;
vram[12'h0d2] = 8'h00;
vram[12'h0d3] = 8'h00;
vram[12'h0d4] = 8'h00;
vram[12'h0d5] = 8'h00;
vram[12'h0d6] = 8'h00;
vram[12'h0d7] = 8'h00;
vram[12'h0d8] = 8'h00;
vram[12'h0d9] = 8'h00;
vram[12'h0da] = 8'h00;
vram[12'h0db] = 8'h00;
vram[12'h0dc] = 8'h00;
vram[12'h0dd] = 8'h00;
vram[12'h0de] = 8'h00;
vram[12'h0df] = 8'h00;
vram[12'h0e0] = 8'h00;
vram[12'h0e1] = 8'h00;
vram[12'h0e2] = 8'h00;
vram[12'h0e3] = 8'h00;
vram[12'h0e4] = 8'h00;
vram[12'h0e5] = 8'h00;
vram[12'h0e6] = 8'h00;
vram[12'h0e7] = 8'h00;
vram[12'h0e8] = 8'h00;
vram[12'h0e9] = 8'h00;
vram[12'h0ea] = 8'h00;
vram[12'h0eb] = 8'h00;
vram[12'h0ec] = 8'h00;
vram[12'h0ed] = 8'h00;
vram[12'h0ee] = 8'h00;
vram[12'h0ef] = 8'h00;
vram[12'h0f0] = 8'h00;
vram[12'h0f1] = 8'h00;
vram[12'h0f2] = 8'h00;
vram[12'h0f3] = 8'h00;
vram[12'h0f4] = 8'h00;
vram[12'h0f5] = 8'h00;
vram[12'h0f6] = 8'h00;
vram[12'h0f7] = 8'h00;
vram[12'h0f8] = 8'h00;
vram[12'h0f9] = 8'h00;
vram[12'h0fa] = 8'h00;
vram[12'h0fb] = 8'h00;
vram[12'h0fc] = 8'h00;
vram[12'h0fd] = 8'h00;
vram[12'h0fe] = 8'h00;
vram[12'h0ff] = 8'h00;
vram[12'h100] = 8'h00;
vram[12'h101] = 8'h00;
vram[12'h102] = 8'h00;
vram[12'h103] = 8'h00;
vram[12'h104] = 8'h00;
vram[12'h105] = 8'h00;
vram[12'h106] = 8'h00;
vram[12'h107] = 8'h00;
vram[12'h108] = 8'h00;
vram[12'h109] = 8'h00;
vram[12'h10a] = 8'h00;
vram[12'h10b] = 8'h00;
vram[12'h10c] = 8'h00;
vram[12'h10d] = 8'h00;
vram[12'h10e] = 8'h00;
vram[12'h10f] = 8'h00;
vram[12'h110] = 8'h00;
vram[12'h111] = 8'h00;
vram[12'h112] = 8'h00;
vram[12'h113] = 8'h00;
vram[12'h114] = 8'h00;
vram[12'h115] = 8'h00;
vram[12'h116] = 8'h00;
vram[12'h117] = 8'h00;
vram[12'h118] = 8'h00;
vram[12'h119] = 8'h00;
vram[12'h11a] = 8'h00;
vram[12'h11b] = 8'h00;
vram[12'h11c] = 8'h00;
vram[12'h11d] = 8'h00;
vram[12'h11e] = 8'h00;
vram[12'h11f] = 8'h00;
vram[12'h120] = 8'h00;
vram[12'h121] = 8'h00;
vram[12'h122] = 8'h00;
vram[12'h123] = 8'h00;
vram[12'h124] = 8'h00;
vram[12'h125] = 8'h00;
vram[12'h126] = 8'h00;
vram[12'h127] = 8'h00;
vram[12'h128] = 8'h00;
vram[12'h129] = 8'h00;
vram[12'h12a] = 8'h00;
vram[12'h12b] = 8'h00;
vram[12'h12c] = 8'h00;
vram[12'h12d] = 8'h00;
vram[12'h12e] = 8'h00;
vram[12'h12f] = 8'h00;
vram[12'h130] = 8'h00;
vram[12'h131] = 8'h00;
vram[12'h132] = 8'h00;
vram[12'h133] = 8'h00;
vram[12'h134] = 8'h00;
vram[12'h135] = 8'h00;
vram[12'h136] = 8'h00;
vram[12'h137] = 8'h00;
vram[12'h138] = 8'h00;
vram[12'h139] = 8'h00;
vram[12'h13a] = 8'h00;
vram[12'h13b] = 8'h00;
vram[12'h13c] = 8'h00;
vram[12'h13d] = 8'h00;
vram[12'h13e] = 8'h00;
vram[12'h13f] = 8'h00;
vram[12'h140] = 8'h00;
vram[12'h141] = 8'h00;
vram[12'h142] = 8'h00;
vram[12'h143] = 8'h00;
vram[12'h144] = 8'h00;
vram[12'h145] = 8'h00;
vram[12'h146] = 8'h00;
vram[12'h147] = 8'h00;
vram[12'h148] = 8'h00;
vram[12'h149] = 8'h00;
vram[12'h14a] = 8'h00;
vram[12'h14b] = 8'h00;
vram[12'h14c] = 8'h00;
vram[12'h14d] = 8'h00;
vram[12'h14e] = 8'h00;
vram[12'h14f] = 8'h00;
vram[12'h150] = 8'h00;
vram[12'h151] = 8'h00;
vram[12'h152] = 8'h00;
vram[12'h153] = 8'h00;
vram[12'h154] = 8'h00;
vram[12'h155] = 8'h00;
vram[12'h156] = 8'h00;
vram[12'h157] = 8'h00;
vram[12'h158] = 8'h00;
vram[12'h159] = 8'h00;
vram[12'h15a] = 8'h00;
vram[12'h15b] = 8'h00;
vram[12'h15c] = 8'h00;
vram[12'h15d] = 8'h00;
vram[12'h15e] = 8'h00;
vram[12'h15f] = 8'h00;
vram[12'h160] = 8'h00;
vram[12'h161] = 8'h00;
vram[12'h162] = 8'h00;
vram[12'h163] = 8'h00;
vram[12'h164] = 8'h00;
vram[12'h165] = 8'h00;
vram[12'h166] = 8'h00;
vram[12'h167] = 8'h00;
vram[12'h168] = 8'h00;
vram[12'h169] = 8'h00;
vram[12'h16a] = 8'h00;
vram[12'h16b] = 8'h00;
vram[12'h16c] = 8'h00;
vram[12'h16d] = 8'h00;
vram[12'h16e] = 8'h00;
vram[12'h16f] = 8'h00;
vram[12'h170] = 8'h00;
vram[12'h171] = 8'h00;
vram[12'h172] = 8'h00;
vram[12'h173] = 8'h00;
vram[12'h174] = 8'h00;
vram[12'h175] = 8'h00;
vram[12'h176] = 8'h00;
vram[12'h177] = 8'h00;
vram[12'h178] = 8'h00;
vram[12'h179] = 8'h00;
vram[12'h17a] = 8'h00;
vram[12'h17b] = 8'h00;
vram[12'h17c] = 8'h00;
vram[12'h17d] = 8'h00;
vram[12'h17e] = 8'h00;
vram[12'h17f] = 8'h00;
vram[12'h180] = 8'h00;
vram[12'h181] = 8'h00;
vram[12'h182] = 8'h00;
vram[12'h183] = 8'h00;
vram[12'h184] = 8'h00;
vram[12'h185] = 8'h00;
vram[12'h186] = 8'h00;
vram[12'h187] = 8'h00;
vram[12'h188] = 8'h00;
vram[12'h189] = 8'h00;
vram[12'h18a] = 8'h00;
vram[12'h18b] = 8'h00;
vram[12'h18c] = 8'h00;
vram[12'h18d] = 8'h00;
vram[12'h18e] = 8'h00;
vram[12'h18f] = 8'h00;
vram[12'h190] = 8'h00;
vram[12'h191] = 8'h00;
vram[12'h192] = 8'h00;
vram[12'h193] = 8'h00;
vram[12'h194] = 8'h00;
vram[12'h195] = 8'h00;
vram[12'h196] = 8'h00;
vram[12'h197] = 8'h00;
vram[12'h198] = 8'h00;
vram[12'h199] = 8'h00;
vram[12'h19a] = 8'h00;
vram[12'h19b] = 8'h00;
vram[12'h19c] = 8'h00;
vram[12'h19d] = 8'h00;
vram[12'h19e] = 8'h00;
vram[12'h19f] = 8'h00;
vram[12'h1a0] = 8'h00;
vram[12'h1a1] = 8'h00;
vram[12'h1a2] = 8'h00;
vram[12'h1a3] = 8'h00;
vram[12'h1a4] = 8'h00;
vram[12'h1a5] = 8'h00;
vram[12'h1a6] = 8'h00;
vram[12'h1a7] = 8'h00;
vram[12'h1a8] = 8'h00;
vram[12'h1a9] = 8'h00;
vram[12'h1aa] = 8'h00;
vram[12'h1ab] = 8'h00;
vram[12'h1ac] = 8'h00;
vram[12'h1ad] = 8'h00;
vram[12'h1ae] = 8'h00;
vram[12'h1af] = 8'h00;
vram[12'h1b0] = 8'h00;
vram[12'h1b1] = 8'h00;
vram[12'h1b2] = 8'h00;
vram[12'h1b3] = 8'h00;
vram[12'h1b4] = 8'h00;
vram[12'h1b5] = 8'h00;
vram[12'h1b6] = 8'h00;
vram[12'h1b7] = 8'h00;
vram[12'h1b8] = 8'h00;
vram[12'h1b9] = 8'h00;
vram[12'h1ba] = 8'h00;
vram[12'h1bb] = 8'h00;
vram[12'h1bc] = 8'h00;
vram[12'h1bd] = 8'h00;
vram[12'h1be] = 8'h00;
vram[12'h1bf] = 8'h00;
vram[12'h1c0] = 8'h00;
vram[12'h1c1] = 8'h00;
vram[12'h1c2] = 8'h00;
vram[12'h1c3] = 8'h00;
vram[12'h1c4] = 8'h00;
vram[12'h1c5] = 8'h00;
vram[12'h1c6] = 8'h00;
vram[12'h1c7] = 8'h00;
vram[12'h1c8] = 8'h00;
vram[12'h1c9] = 8'h00;
vram[12'h1ca] = 8'h00;
vram[12'h1cb] = 8'h00;
vram[12'h1cc] = 8'h00;
vram[12'h1cd] = 8'h00;
vram[12'h1ce] = 8'h00;
vram[12'h1cf] = 8'h00;
vram[12'h1d0] = 8'h00;
vram[12'h1d1] = 8'h00;
vram[12'h1d2] = 8'h00;
vram[12'h1d3] = 8'h00;
vram[12'h1d4] = 8'h00;
vram[12'h1d5] = 8'h00;
vram[12'h1d6] = 8'h00;
vram[12'h1d7] = 8'h00;
vram[12'h1d8] = 8'h00;
vram[12'h1d9] = 8'h00;
vram[12'h1da] = 8'h00;
vram[12'h1db] = 8'h00;
vram[12'h1dc] = 8'h00;
vram[12'h1dd] = 8'h00;
vram[12'h1de] = 8'h00;
vram[12'h1df] = 8'h00;
vram[12'h1e0] = 8'h00;
vram[12'h1e1] = 8'h00;
vram[12'h1e2] = 8'h00;
vram[12'h1e3] = 8'h00;
vram[12'h1e4] = 8'h00;
vram[12'h1e5] = 8'h00;
vram[12'h1e6] = 8'h00;
vram[12'h1e7] = 8'h00;
vram[12'h1e8] = 8'h00;
vram[12'h1e9] = 8'h00;
vram[12'h1ea] = 8'h00;
vram[12'h1eb] = 8'h00;
vram[12'h1ec] = 8'h00;
vram[12'h1ed] = 8'h00;
vram[12'h1ee] = 8'h00;
vram[12'h1ef] = 8'h00;
vram[12'h1f0] = 8'h00;
vram[12'h1f1] = 8'h00;
vram[12'h1f2] = 8'h00;
vram[12'h1f3] = 8'h00;
vram[12'h1f4] = 8'h00;
vram[12'h1f5] = 8'h00;
vram[12'h1f6] = 8'h00;
vram[12'h1f7] = 8'h00;
vram[12'h1f8] = 8'h00;
vram[12'h1f9] = 8'h00;
vram[12'h1fa] = 8'h00;
vram[12'h1fb] = 8'h00;
vram[12'h1fc] = 8'h00;
vram[12'h1fd] = 8'h00;
vram[12'h1fe] = 8'h00;
vram[12'h1ff] = 8'h00;
vram[12'h200] = 8'h00;
vram[12'h201] = 8'h00;
vram[12'h202] = 8'h00;
vram[12'h203] = 8'h00;
vram[12'h204] = 8'h00;
vram[12'h205] = 8'h00;
vram[12'h206] = 8'h00;
vram[12'h207] = 8'h00;
vram[12'h208] = 8'h00;
vram[12'h209] = 8'h00;
vram[12'h20a] = 8'h00;
vram[12'h20b] = 8'h00;
vram[12'h20c] = 8'h00;
vram[12'h20d] = 8'h00;
vram[12'h20e] = 8'h00;
vram[12'h20f] = 8'h00;
vram[12'h210] = 8'h00;
vram[12'h211] = 8'h00;
vram[12'h212] = 8'h00;
vram[12'h213] = 8'h00;
vram[12'h214] = 8'h00;
vram[12'h215] = 8'h00;
vram[12'h216] = 8'h00;
vram[12'h217] = 8'h00;
vram[12'h218] = 8'h00;
vram[12'h219] = 8'h00;
vram[12'h21a] = 8'h00;
vram[12'h21b] = 8'h00;
vram[12'h21c] = 8'h00;
vram[12'h21d] = 8'h00;
vram[12'h21e] = 8'h00;
vram[12'h21f] = 8'h00;
vram[12'h220] = 8'h00;
vram[12'h221] = 8'h00;
vram[12'h222] = 8'h00;
vram[12'h223] = 8'h00;
vram[12'h224] = 8'h00;
vram[12'h225] = 8'h00;
vram[12'h226] = 8'h00;
vram[12'h227] = 8'h00;
vram[12'h228] = 8'h00;
vram[12'h229] = 8'h00;
vram[12'h22a] = 8'h00;
vram[12'h22b] = 8'h00;
vram[12'h22c] = 8'h00;
vram[12'h22d] = 8'h00;
vram[12'h22e] = 8'h00;
vram[12'h22f] = 8'h00;
vram[12'h230] = 8'h00;
vram[12'h231] = 8'h00;
vram[12'h232] = 8'h00;
vram[12'h233] = 8'h00;
vram[12'h234] = 8'h00;
vram[12'h235] = 8'h00;
vram[12'h236] = 8'h00;
vram[12'h237] = 8'h00;
vram[12'h238] = 8'h00;
vram[12'h239] = 8'h00;
vram[12'h23a] = 8'h00;
vram[12'h23b] = 8'h00;
vram[12'h23c] = 8'h00;
vram[12'h23d] = 8'h00;
vram[12'h23e] = 8'h00;
vram[12'h23f] = 8'h00;
vram[12'h240] = 8'h00;
vram[12'h241] = 8'h00;
vram[12'h242] = 8'h00;
vram[12'h243] = 8'h00;
vram[12'h244] = 8'h00;
vram[12'h245] = 8'h00;
vram[12'h246] = 8'h00;
vram[12'h247] = 8'h00;
vram[12'h248] = 8'h00;
vram[12'h249] = 8'h00;
vram[12'h24a] = 8'h00;
vram[12'h24b] = 8'h00;
vram[12'h24c] = 8'h00;
vram[12'h24d] = 8'h00;
vram[12'h24e] = 8'h00;
vram[12'h24f] = 8'h00;
vram[12'h250] = 8'h00;
vram[12'h251] = 8'h00;
vram[12'h252] = 8'h00;
vram[12'h253] = 8'h00;
vram[12'h254] = 8'h00;
vram[12'h255] = 8'h00;
vram[12'h256] = 8'h00;
vram[12'h257] = 8'h00;
vram[12'h258] = 8'h00;
vram[12'h259] = 8'h00;
vram[12'h25a] = 8'h00;
vram[12'h25b] = 8'h00;
vram[12'h25c] = 8'h00;
vram[12'h25d] = 8'h00;
vram[12'h25e] = 8'h00;
vram[12'h25f] = 8'h00;
vram[12'h260] = 8'h00;
vram[12'h261] = 8'h00;
vram[12'h262] = 8'h00;
vram[12'h263] = 8'h00;
vram[12'h264] = 8'h00;
vram[12'h265] = 8'h00;
vram[12'h266] = 8'h00;
vram[12'h267] = 8'h00;
vram[12'h268] = 8'h00;
vram[12'h269] = 8'h00;
vram[12'h26a] = 8'h00;
vram[12'h26b] = 8'h00;
vram[12'h26c] = 8'h00;
vram[12'h26d] = 8'h00;
vram[12'h26e] = 8'h00;
vram[12'h26f] = 8'h00;
vram[12'h270] = 8'h00;
vram[12'h271] = 8'h00;
vram[12'h272] = 8'h00;
vram[12'h273] = 8'h00;
vram[12'h274] = 8'h00;
vram[12'h275] = 8'h00;
vram[12'h276] = 8'h00;
vram[12'h277] = 8'h00;
vram[12'h278] = 8'h00;
vram[12'h279] = 8'h00;
vram[12'h27a] = 8'h00;
vram[12'h27b] = 8'h00;
vram[12'h27c] = 8'h00;
vram[12'h27d] = 8'h00;
vram[12'h27e] = 8'h00;
vram[12'h27f] = 8'h00;
vram[12'h280] = 8'h00;
vram[12'h281] = 8'h00;
vram[12'h282] = 8'h00;
vram[12'h283] = 8'h00;
vram[12'h284] = 8'h00;
vram[12'h285] = 8'h00;
vram[12'h286] = 8'h00;
vram[12'h287] = 8'h00;
vram[12'h288] = 8'h00;
vram[12'h289] = 8'h00;
vram[12'h28a] = 8'h00;
vram[12'h28b] = 8'h00;
vram[12'h28c] = 8'h00;
vram[12'h28d] = 8'h00;
vram[12'h28e] = 8'h00;
vram[12'h28f] = 8'h00;
vram[12'h290] = 8'h00;
vram[12'h291] = 8'h00;
vram[12'h292] = 8'h00;
vram[12'h293] = 8'h00;
vram[12'h294] = 8'h00;
vram[12'h295] = 8'h00;
vram[12'h296] = 8'h00;
vram[12'h297] = 8'h00;
vram[12'h298] = 8'h00;
vram[12'h299] = 8'h00;
vram[12'h29a] = 8'h00;
vram[12'h29b] = 8'h00;
vram[12'h29c] = 8'h00;
vram[12'h29d] = 8'h00;
vram[12'h29e] = 8'h00;
vram[12'h29f] = 8'h00;
vram[12'h2a0] = 8'h00;
vram[12'h2a1] = 8'h00;
vram[12'h2a2] = 8'h00;
vram[12'h2a3] = 8'h00;
vram[12'h2a4] = 8'h00;
vram[12'h2a5] = 8'h00;
vram[12'h2a6] = 8'h00;
vram[12'h2a7] = 8'h00;
vram[12'h2a8] = 8'h00;
vram[12'h2a9] = 8'h00;
vram[12'h2aa] = 8'h00;
vram[12'h2ab] = 8'h00;
vram[12'h2ac] = 8'h00;
vram[12'h2ad] = 8'h00;
vram[12'h2ae] = 8'h00;
vram[12'h2af] = 8'h00;
vram[12'h2b0] = 8'h00;
vram[12'h2b1] = 8'h00;
vram[12'h2b2] = 8'h00;
vram[12'h2b3] = 8'h00;
vram[12'h2b4] = 8'h00;
vram[12'h2b5] = 8'h00;
vram[12'h2b6] = 8'h00;
vram[12'h2b7] = 8'h00;
vram[12'h2b8] = 8'h00;
vram[12'h2b9] = 8'h00;
vram[12'h2ba] = 8'h00;
vram[12'h2bb] = 8'h00;
vram[12'h2bc] = 8'h00;
vram[12'h2bd] = 8'h00;
vram[12'h2be] = 8'h00;
vram[12'h2bf] = 8'h00;
vram[12'h2c0] = 8'h00;
vram[12'h2c1] = 8'h00;
vram[12'h2c2] = 8'h00;
vram[12'h2c3] = 8'h00;
vram[12'h2c4] = 8'h00;
vram[12'h2c5] = 8'h00;
vram[12'h2c6] = 8'h00;
vram[12'h2c7] = 8'h00;
vram[12'h2c8] = 8'h00;
vram[12'h2c9] = 8'h00;
vram[12'h2ca] = 8'h00;
vram[12'h2cb] = 8'h00;
vram[12'h2cc] = 8'h00;
vram[12'h2cd] = 8'h00;
vram[12'h2ce] = 8'h00;
vram[12'h2cf] = 8'h00;
vram[12'h2d0] = 8'h00;
vram[12'h2d1] = 8'h00;
vram[12'h2d2] = 8'h00;
vram[12'h2d3] = 8'h00;
vram[12'h2d4] = 8'h00;
vram[12'h2d5] = 8'h00;
vram[12'h2d6] = 8'h00;
vram[12'h2d7] = 8'h00;
vram[12'h2d8] = 8'h00;
vram[12'h2d9] = 8'h00;
vram[12'h2da] = 8'h00;
vram[12'h2db] = 8'h00;
vram[12'h2dc] = 8'h00;
vram[12'h2dd] = 8'h00;
vram[12'h2de] = 8'h00;
vram[12'h2df] = 8'h00;
vram[12'h2e0] = 8'h00;
vram[12'h2e1] = 8'h00;
vram[12'h2e2] = 8'h00;
vram[12'h2e3] = 8'h00;
vram[12'h2e4] = 8'h00;
vram[12'h2e5] = 8'h00;
vram[12'h2e6] = 8'h00;
vram[12'h2e7] = 8'h00;
vram[12'h2e8] = 8'h00;
vram[12'h2e9] = 8'h00;
vram[12'h2ea] = 8'h00;
vram[12'h2eb] = 8'h00;
vram[12'h2ec] = 8'h00;
vram[12'h2ed] = 8'h00;
vram[12'h2ee] = 8'h00;
vram[12'h2ef] = 8'h00;
vram[12'h2f0] = 8'h00;
vram[12'h2f1] = 8'h00;
vram[12'h2f2] = 8'h00;
vram[12'h2f3] = 8'h00;
vram[12'h2f4] = 8'h00;
vram[12'h2f5] = 8'h00;
vram[12'h2f6] = 8'h00;
vram[12'h2f7] = 8'h00;
vram[12'h2f8] = 8'h00;
vram[12'h2f9] = 8'h00;
vram[12'h2fa] = 8'h00;
vram[12'h2fb] = 8'h00;
vram[12'h2fc] = 8'h00;
vram[12'h2fd] = 8'h00;
vram[12'h2fe] = 8'h00;
vram[12'h2ff] = 8'h00;
vram[12'h300] = 8'h00;
vram[12'h301] = 8'h00;
vram[12'h302] = 8'h00;
vram[12'h303] = 8'h00;
vram[12'h304] = 8'h00;
vram[12'h305] = 8'h00;
vram[12'h306] = 8'h00;
vram[12'h307] = 8'h00;
vram[12'h308] = 8'h00;
vram[12'h309] = 8'h00;
vram[12'h30a] = 8'h00;
vram[12'h30b] = 8'h00;
vram[12'h30c] = 8'h00;
vram[12'h30d] = 8'h00;
vram[12'h30e] = 8'h00;
vram[12'h30f] = 8'h00;
vram[12'h310] = 8'h00;
vram[12'h311] = 8'h00;
vram[12'h312] = 8'h00;
vram[12'h313] = 8'h00;
vram[12'h314] = 8'h00;
vram[12'h315] = 8'h00;
vram[12'h316] = 8'h00;
vram[12'h317] = 8'h00;
vram[12'h318] = 8'h00;
vram[12'h319] = 8'h00;
vram[12'h31a] = 8'h00;
vram[12'h31b] = 8'h00;
vram[12'h31c] = 8'h00;
vram[12'h31d] = 8'h00;
vram[12'h31e] = 8'h00;
vram[12'h31f] = 8'h00;
vram[12'h320] = 8'h00;
vram[12'h321] = 8'h00;
vram[12'h322] = 8'h00;
vram[12'h323] = 8'h00;
vram[12'h324] = 8'h00;
vram[12'h325] = 8'h00;
vram[12'h326] = 8'h00;
vram[12'h327] = 8'h00;
vram[12'h328] = 8'h00;
vram[12'h329] = 8'h00;
vram[12'h32a] = 8'h00;
vram[12'h32b] = 8'h00;
vram[12'h32c] = 8'h00;
vram[12'h32d] = 8'h00;
vram[12'h32e] = 8'h00;
vram[12'h32f] = 8'h00;
vram[12'h330] = 8'h00;
vram[12'h331] = 8'h00;
vram[12'h332] = 8'h00;
vram[12'h333] = 8'h00;
vram[12'h334] = 8'h00;
vram[12'h335] = 8'h00;
vram[12'h336] = 8'h00;
vram[12'h337] = 8'h00;
vram[12'h338] = 8'h00;
vram[12'h339] = 8'h00;
vram[12'h33a] = 8'h00;
vram[12'h33b] = 8'h00;
vram[12'h33c] = 8'h00;
vram[12'h33d] = 8'h00;
vram[12'h33e] = 8'h00;
vram[12'h33f] = 8'h00;
vram[12'h340] = 8'h00;
vram[12'h341] = 8'h00;
vram[12'h342] = 8'h00;
vram[12'h343] = 8'h00;
vram[12'h344] = 8'h00;
vram[12'h345] = 8'h00;
vram[12'h346] = 8'h00;
vram[12'h347] = 8'h00;
vram[12'h348] = 8'h00;
vram[12'h349] = 8'h00;
vram[12'h34a] = 8'h00;
vram[12'h34b] = 8'h00;
vram[12'h34c] = 8'h00;
vram[12'h34d] = 8'h00;
vram[12'h34e] = 8'h00;
vram[12'h34f] = 8'h00;
vram[12'h350] = 8'h00;
vram[12'h351] = 8'h00;
vram[12'h352] = 8'h00;
vram[12'h353] = 8'h00;
vram[12'h354] = 8'h00;
vram[12'h355] = 8'h00;
vram[12'h356] = 8'h00;
vram[12'h357] = 8'h00;
vram[12'h358] = 8'h00;
vram[12'h359] = 8'h00;
vram[12'h35a] = 8'h00;
vram[12'h35b] = 8'h00;
vram[12'h35c] = 8'h00;
vram[12'h35d] = 8'h00;
vram[12'h35e] = 8'h00;
vram[12'h35f] = 8'h00;
vram[12'h360] = 8'h00;
vram[12'h361] = 8'h00;
vram[12'h362] = 8'h00;
vram[12'h363] = 8'h00;
vram[12'h364] = 8'h00;
vram[12'h365] = 8'h00;
vram[12'h366] = 8'h00;
vram[12'h367] = 8'h00;
vram[12'h368] = 8'h00;
vram[12'h369] = 8'h00;
vram[12'h36a] = 8'h00;
vram[12'h36b] = 8'h00;
vram[12'h36c] = 8'h00;
vram[12'h36d] = 8'h00;
vram[12'h36e] = 8'h00;
vram[12'h36f] = 8'h00;
vram[12'h370] = 8'h00;
vram[12'h371] = 8'h00;
vram[12'h372] = 8'h00;
vram[12'h373] = 8'h00;
vram[12'h374] = 8'h00;
vram[12'h375] = 8'h00;
vram[12'h376] = 8'h00;
vram[12'h377] = 8'h00;
vram[12'h378] = 8'h00;
vram[12'h379] = 8'h00;
vram[12'h37a] = 8'h00;
vram[12'h37b] = 8'h00;
vram[12'h37c] = 8'h00;
vram[12'h37d] = 8'h00;
vram[12'h37e] = 8'h00;
vram[12'h37f] = 8'h00;
vram[12'h380] = 8'h00;
vram[12'h381] = 8'h00;
vram[12'h382] = 8'h00;
vram[12'h383] = 8'h00;
vram[12'h384] = 8'h00;
vram[12'h385] = 8'h00;
vram[12'h386] = 8'h00;
vram[12'h387] = 8'h00;
vram[12'h388] = 8'h00;
vram[12'h389] = 8'h00;
vram[12'h38a] = 8'h00;
vram[12'h38b] = 8'h00;
vram[12'h38c] = 8'h00;
vram[12'h38d] = 8'h00;
vram[12'h38e] = 8'h00;
vram[12'h38f] = 8'h00;
vram[12'h390] = 8'h00;
vram[12'h391] = 8'h00;
vram[12'h392] = 8'h00;
vram[12'h393] = 8'h00;
vram[12'h394] = 8'h00;
vram[12'h395] = 8'h00;
vram[12'h396] = 8'h00;
vram[12'h397] = 8'h00;
vram[12'h398] = 8'h00;
vram[12'h399] = 8'h00;
vram[12'h39a] = 8'h00;
vram[12'h39b] = 8'h00;
vram[12'h39c] = 8'h00;
vram[12'h39d] = 8'h00;
vram[12'h39e] = 8'h00;
vram[12'h39f] = 8'h00;
vram[12'h3a0] = 8'h00;
vram[12'h3a1] = 8'h00;
vram[12'h3a2] = 8'h00;
vram[12'h3a3] = 8'h00;
vram[12'h3a4] = 8'h00;
vram[12'h3a5] = 8'h00;
vram[12'h3a6] = 8'h00;
vram[12'h3a7] = 8'h00;
vram[12'h3a8] = 8'h00;
vram[12'h3a9] = 8'h00;
vram[12'h3aa] = 8'h00;
vram[12'h3ab] = 8'h00;
vram[12'h3ac] = 8'h00;
vram[12'h3ad] = 8'h00;
vram[12'h3ae] = 8'h00;
vram[12'h3af] = 8'h00;
vram[12'h3b0] = 8'h00;
vram[12'h3b1] = 8'h00;
vram[12'h3b2] = 8'h00;
vram[12'h3b3] = 8'h00;
vram[12'h3b4] = 8'h00;
vram[12'h3b5] = 8'h00;
vram[12'h3b6] = 8'h00;
vram[12'h3b7] = 8'h00;
vram[12'h3b8] = 8'h00;
vram[12'h3b9] = 8'h00;
vram[12'h3ba] = 8'h00;
vram[12'h3bb] = 8'h00;
vram[12'h3bc] = 8'h00;
vram[12'h3bd] = 8'h00;
vram[12'h3be] = 8'h00;
vram[12'h3bf] = 8'h00;
vram[12'h3c0] = 8'h00;
vram[12'h3c1] = 8'h00;
vram[12'h3c2] = 8'h00;
vram[12'h3c3] = 8'h00;
vram[12'h3c4] = 8'h00;
vram[12'h3c5] = 8'h00;
vram[12'h3c6] = 8'h00;
vram[12'h3c7] = 8'h00;
vram[12'h3c8] = 8'h00;
vram[12'h3c9] = 8'h00;
vram[12'h3ca] = 8'h00;
vram[12'h3cb] = 8'h00;
vram[12'h3cc] = 8'h00;
vram[12'h3cd] = 8'h00;
vram[12'h3ce] = 8'h00;
vram[12'h3cf] = 8'h00;
vram[12'h3d0] = 8'h00;
vram[12'h3d1] = 8'h00;
vram[12'h3d2] = 8'h00;
vram[12'h3d3] = 8'h00;
vram[12'h3d4] = 8'h00;
vram[12'h3d5] = 8'h00;
vram[12'h3d6] = 8'h00;
vram[12'h3d7] = 8'h00;
vram[12'h3d8] = 8'h00;
vram[12'h3d9] = 8'h00;
vram[12'h3da] = 8'h00;
vram[12'h3db] = 8'h00;
vram[12'h3dc] = 8'h00;
vram[12'h3dd] = 8'h00;
vram[12'h3de] = 8'h00;
vram[12'h3df] = 8'h00;
vram[12'h3e0] = 8'h00;
vram[12'h3e1] = 8'h00;
vram[12'h3e2] = 8'h00;
vram[12'h3e3] = 8'h00;
vram[12'h3e4] = 8'h00;
vram[12'h3e5] = 8'h00;
vram[12'h3e6] = 8'h00;
vram[12'h3e7] = 8'h00;
vram[12'h3e8] = 8'h00;
vram[12'h3e9] = 8'h00;
vram[12'h3ea] = 8'h00;
vram[12'h3eb] = 8'h00;
vram[12'h3ec] = 8'h00;
vram[12'h3ed] = 8'h00;
vram[12'h3ee] = 8'h00;
vram[12'h3ef] = 8'h00;
vram[12'h3f0] = 8'h00;
vram[12'h3f1] = 8'h00;
vram[12'h3f2] = 8'h00;
vram[12'h3f3] = 8'h00;
vram[12'h3f4] = 8'h00;
vram[12'h3f5] = 8'h00;
vram[12'h3f6] = 8'h00;
vram[12'h3f7] = 8'h00;
vram[12'h3f8] = 8'h00;
vram[12'h3f9] = 8'h00;
vram[12'h3fa] = 8'h00;
vram[12'h3fb] = 8'h00;
vram[12'h3fc] = 8'h00;
vram[12'h3fd] = 8'h00;
vram[12'h3fe] = 8'h00;
vram[12'h3ff] = 8'h00;
vram[12'h400] = 8'h00;
vram[12'h401] = 8'h01;
vram[12'h402] = 8'h02;
vram[12'h403] = 8'h03;
vram[12'h404] = 8'h04;
vram[12'h405] = 8'h05;
vram[12'h406] = 8'h06;
vram[12'h407] = 8'h07;
vram[12'h408] = 8'h08;
vram[12'h409] = 8'h09;
vram[12'h40a] = 8'h0a;
vram[12'h40b] = 8'h0b;
vram[12'h40c] = 8'h0c;
vram[12'h40d] = 8'h0d;
vram[12'h40e] = 8'h0e;
vram[12'h40f] = 8'h0f;
vram[12'h410] = 8'h0f;
vram[12'h411] = 8'h0e;
vram[12'h412] = 8'h0d;
vram[12'h413] = 8'h0c;
vram[12'h414] = 8'h0b;
vram[12'h415] = 8'h0a;
vram[12'h416] = 8'h09;
vram[12'h417] = 8'h08;
vram[12'h418] = 8'h07;
vram[12'h419] = 8'h06;
vram[12'h41a] = 8'h05;
vram[12'h41b] = 8'h04;
vram[12'h41c] = 8'h03;
vram[12'h41d] = 8'h02;
vram[12'h41e] = 8'h01;
vram[12'h41f] = 8'h00;
vram[12'h420] = 8'h0f;
vram[12'h421] = 8'h0f;
vram[12'h422] = 8'h0f;
vram[12'h423] = 8'h0f;
vram[12'h424] = 8'h0f;
vram[12'h425] = 8'h0f;
vram[12'h426] = 8'h0f;
vram[12'h427] = 8'h0f;
vram[12'h428] = 8'h0f;
vram[12'h429] = 8'h0f;
vram[12'h42a] = 8'h0f;
vram[12'h42b] = 8'h0f;
vram[12'h42c] = 8'h0f;
vram[12'h42d] = 8'h0f;
vram[12'h42e] = 8'h0f;
vram[12'h42f] = 8'h0f;
vram[12'h430] = 8'h0f;
vram[12'h431] = 8'h0f;
vram[12'h432] = 8'h0f;
vram[12'h433] = 8'h0f;
vram[12'h434] = 8'h0f;
vram[12'h435] = 8'h0f;
vram[12'h436] = 8'h0f;
vram[12'h437] = 8'h0f;
vram[12'h438] = 8'h0f;
vram[12'h439] = 8'h0f;
vram[12'h43a] = 8'h0f;
vram[12'h43b] = 8'h0f;
vram[12'h43c] = 8'h0f;
vram[12'h43d] = 8'h0f;
vram[12'h43e] = 8'h0f;
vram[12'h43f] = 8'h0f;
vram[12'h440] = 8'h0f;
vram[12'h441] = 8'h0f;
vram[12'h442] = 8'h0f;
vram[12'h443] = 8'h0f;
vram[12'h444] = 8'h0f;
vram[12'h445] = 8'h0f;
vram[12'h446] = 8'h0f;
vram[12'h447] = 8'h0f;
vram[12'h448] = 8'h0f;
vram[12'h449] = 8'h0f;
vram[12'h44a] = 8'h0f;
vram[12'h44b] = 8'h0f;
vram[12'h44c] = 8'h0f;
vram[12'h44d] = 8'h0f;
vram[12'h44e] = 8'h0f;
vram[12'h44f] = 8'h0f;
vram[12'h450] = 8'h0f;
vram[12'h451] = 8'h0f;
vram[12'h452] = 8'h0f;
vram[12'h453] = 8'h0f;
vram[12'h454] = 8'h0f;
vram[12'h455] = 8'h0f;
vram[12'h456] = 8'h0f;
vram[12'h457] = 8'h0f;
vram[12'h458] = 8'h0f;
vram[12'h459] = 8'h0f;
vram[12'h45a] = 8'h0f;
vram[12'h45b] = 8'h0f;
vram[12'h45c] = 8'h0f;
vram[12'h45d] = 8'h0f;
vram[12'h45e] = 8'h0f;
vram[12'h45f] = 8'h0f;
vram[12'h460] = 8'h0f;
vram[12'h461] = 8'h0f;
vram[12'h462] = 8'h0f;
vram[12'h463] = 8'h0f;
vram[12'h464] = 8'h0f;
vram[12'h465] = 8'h0f;
vram[12'h466] = 8'h0f;
vram[12'h467] = 8'h0f;
vram[12'h468] = 8'h0f;
vram[12'h469] = 8'h0f;
vram[12'h46a] = 8'h0f;
vram[12'h46b] = 8'h0f;
vram[12'h46c] = 8'h0f;
vram[12'h46d] = 8'h0f;
vram[12'h46e] = 8'h0f;
vram[12'h46f] = 8'h0f;
vram[12'h470] = 8'h0f;
vram[12'h471] = 8'h0f;
vram[12'h472] = 8'h0f;
vram[12'h473] = 8'h0f;
vram[12'h474] = 8'h0f;
vram[12'h475] = 8'h0f;
vram[12'h476] = 8'h0f;
vram[12'h477] = 8'h0f;
vram[12'h478] = 8'h0f;
vram[12'h479] = 8'h0f;
vram[12'h47a] = 8'h0f;
vram[12'h47b] = 8'h0f;
vram[12'h47c] = 8'h0f;
vram[12'h47d] = 8'h0f;
vram[12'h47e] = 8'h0f;
vram[12'h47f] = 8'h0f;
vram[12'h480] = 8'h0f;
vram[12'h481] = 8'h0f;
vram[12'h482] = 8'h0f;
vram[12'h483] = 8'h0f;
vram[12'h484] = 8'h0f;
vram[12'h485] = 8'h0f;
vram[12'h486] = 8'h0f;
vram[12'h487] = 8'h0f;
vram[12'h488] = 8'h0f;
vram[12'h489] = 8'h0f;
vram[12'h48a] = 8'h0f;
vram[12'h48b] = 8'h0f;
vram[12'h48c] = 8'h0f;
vram[12'h48d] = 8'h0f;
vram[12'h48e] = 8'h0f;
vram[12'h48f] = 8'h0f;
vram[12'h490] = 8'h0f;
vram[12'h491] = 8'h0f;
vram[12'h492] = 8'h0f;
vram[12'h493] = 8'h0f;
vram[12'h494] = 8'h0f;
vram[12'h495] = 8'h0f;
vram[12'h496] = 8'h0f;
vram[12'h497] = 8'h0f;
vram[12'h498] = 8'h0f;
vram[12'h499] = 8'h0f;
vram[12'h49a] = 8'h0f;
vram[12'h49b] = 8'h0f;
vram[12'h49c] = 8'h0f;
vram[12'h49d] = 8'h0f;
vram[12'h49e] = 8'h0f;
vram[12'h49f] = 8'h0f;
vram[12'h4a0] = 8'h0f;
vram[12'h4a1] = 8'h0f;
vram[12'h4a2] = 8'h0f;
vram[12'h4a3] = 8'h0f;
vram[12'h4a4] = 8'h0f;
vram[12'h4a5] = 8'h0f;
vram[12'h4a6] = 8'h0f;
vram[12'h4a7] = 8'h0f;
vram[12'h4a8] = 8'h0f;
vram[12'h4a9] = 8'h0f;
vram[12'h4aa] = 8'h0f;
vram[12'h4ab] = 8'h0f;
vram[12'h4ac] = 8'h0f;
vram[12'h4ad] = 8'h0f;
vram[12'h4ae] = 8'h0f;
vram[12'h4af] = 8'h0f;
vram[12'h4b0] = 8'h0f;
vram[12'h4b1] = 8'h0f;
vram[12'h4b2] = 8'h0f;
vram[12'h4b3] = 8'h0f;
vram[12'h4b4] = 8'h0f;
vram[12'h4b5] = 8'h0f;
vram[12'h4b6] = 8'h0f;
vram[12'h4b7] = 8'h0f;
vram[12'h4b8] = 8'h0f;
vram[12'h4b9] = 8'h0f;
vram[12'h4ba] = 8'h0f;
vram[12'h4bb] = 8'h0f;
vram[12'h4bc] = 8'h0f;
vram[12'h4bd] = 8'h0f;
vram[12'h4be] = 8'h0f;
vram[12'h4bf] = 8'h0f;
vram[12'h4c0] = 8'h0f;
vram[12'h4c1] = 8'h0f;
vram[12'h4c2] = 8'h0f;
vram[12'h4c3] = 8'h0f;
vram[12'h4c4] = 8'h0f;
vram[12'h4c5] = 8'h0f;
vram[12'h4c6] = 8'h0f;
vram[12'h4c7] = 8'h0f;
vram[12'h4c8] = 8'h0f;
vram[12'h4c9] = 8'h0f;
vram[12'h4ca] = 8'h0f;
vram[12'h4cb] = 8'h0f;
vram[12'h4cc] = 8'h0f;
vram[12'h4cd] = 8'h0f;
vram[12'h4ce] = 8'h0f;
vram[12'h4cf] = 8'h0f;
vram[12'h4d0] = 8'h0f;
vram[12'h4d1] = 8'h0f;
vram[12'h4d2] = 8'h0f;
vram[12'h4d3] = 8'h0f;
vram[12'h4d4] = 8'h0f;
vram[12'h4d5] = 8'h0f;
vram[12'h4d6] = 8'h0f;
vram[12'h4d7] = 8'h0f;
vram[12'h4d8] = 8'h0f;
vram[12'h4d9] = 8'h0f;
vram[12'h4da] = 8'h0f;
vram[12'h4db] = 8'h0f;
vram[12'h4dc] = 8'h0f;
vram[12'h4dd] = 8'h0f;
vram[12'h4de] = 8'h0f;
vram[12'h4df] = 8'h0f;
vram[12'h4e0] = 8'h0f;
vram[12'h4e1] = 8'h0f;
vram[12'h4e2] = 8'h0f;
vram[12'h4e3] = 8'h0f;
vram[12'h4e4] = 8'h0f;
vram[12'h4e5] = 8'h0f;
vram[12'h4e6] = 8'h0f;
vram[12'h4e7] = 8'h0f;
vram[12'h4e8] = 8'h0f;
vram[12'h4e9] = 8'h0f;
vram[12'h4ea] = 8'h0f;
vram[12'h4eb] = 8'h0f;
vram[12'h4ec] = 8'h0f;
vram[12'h4ed] = 8'h0f;
vram[12'h4ee] = 8'h0f;
vram[12'h4ef] = 8'h0f;
vram[12'h4f0] = 8'h0f;
vram[12'h4f1] = 8'h0f;
vram[12'h4f2] = 8'h0f;
vram[12'h4f3] = 8'h0f;
vram[12'h4f4] = 8'h0f;
vram[12'h4f5] = 8'h0f;
vram[12'h4f6] = 8'h0f;
vram[12'h4f7] = 8'h0f;
vram[12'h4f8] = 8'h0f;
vram[12'h4f9] = 8'h0f;
vram[12'h4fa] = 8'h0f;
vram[12'h4fb] = 8'h0f;
vram[12'h4fc] = 8'h0f;
vram[12'h4fd] = 8'h0f;
vram[12'h4fe] = 8'h0f;
vram[12'h4ff] = 8'h0f;
vram[12'h500] = 8'h0f;
vram[12'h501] = 8'h0f;
vram[12'h502] = 8'h0f;
vram[12'h503] = 8'h0f;
vram[12'h504] = 8'h0f;
vram[12'h505] = 8'h0f;
vram[12'h506] = 8'h0f;
vram[12'h507] = 8'h0f;
vram[12'h508] = 8'h0f;
vram[12'h509] = 8'h0f;
vram[12'h50a] = 8'h0f;
vram[12'h50b] = 8'h0f;
vram[12'h50c] = 8'h0f;
vram[12'h50d] = 8'h0f;
vram[12'h50e] = 8'h0f;
vram[12'h50f] = 8'h0f;
vram[12'h510] = 8'h0f;
vram[12'h511] = 8'h0f;
vram[12'h512] = 8'h0f;
vram[12'h513] = 8'h0f;
vram[12'h514] = 8'h0f;
vram[12'h515] = 8'h0f;
vram[12'h516] = 8'h0f;
vram[12'h517] = 8'h0f;
vram[12'h518] = 8'h0f;
vram[12'h519] = 8'h0f;
vram[12'h51a] = 8'h0f;
vram[12'h51b] = 8'h0f;
vram[12'h51c] = 8'h0f;
vram[12'h51d] = 8'h0f;
vram[12'h51e] = 8'h0f;
vram[12'h51f] = 8'h0f;
vram[12'h520] = 8'h0f;
vram[12'h521] = 8'h0f;
vram[12'h522] = 8'h0f;
vram[12'h523] = 8'h0f;
vram[12'h524] = 8'h0f;
vram[12'h525] = 8'h0f;
vram[12'h526] = 8'h0f;
vram[12'h527] = 8'h0f;
vram[12'h528] = 8'h0f;
vram[12'h529] = 8'h0f;
vram[12'h52a] = 8'h0f;
vram[12'h52b] = 8'h0f;
vram[12'h52c] = 8'h0f;
vram[12'h52d] = 8'h0f;
vram[12'h52e] = 8'h0f;
vram[12'h52f] = 8'h0f;
vram[12'h530] = 8'h0f;
vram[12'h531] = 8'h0f;
vram[12'h532] = 8'h0f;
vram[12'h533] = 8'h0f;
vram[12'h534] = 8'h0f;
vram[12'h535] = 8'h0f;
vram[12'h536] = 8'h0f;
vram[12'h537] = 8'h0f;
vram[12'h538] = 8'h0f;
vram[12'h539] = 8'h0f;
vram[12'h53a] = 8'h0f;
vram[12'h53b] = 8'h0f;
vram[12'h53c] = 8'h0f;
vram[12'h53d] = 8'h0f;
vram[12'h53e] = 8'h0f;
vram[12'h53f] = 8'h0f;
vram[12'h540] = 8'h0f;
vram[12'h541] = 8'h0f;
vram[12'h542] = 8'h0f;
vram[12'h543] = 8'h0f;
vram[12'h544] = 8'h0f;
vram[12'h545] = 8'h0f;
vram[12'h546] = 8'h0f;
vram[12'h547] = 8'h0f;
vram[12'h548] = 8'h0f;
vram[12'h549] = 8'h0f;
vram[12'h54a] = 8'h0f;
vram[12'h54b] = 8'h0f;
vram[12'h54c] = 8'h0f;
vram[12'h54d] = 8'h0f;
vram[12'h54e] = 8'h0f;
vram[12'h54f] = 8'h0f;
vram[12'h550] = 8'h0f;
vram[12'h551] = 8'h0f;
vram[12'h552] = 8'h0f;
vram[12'h553] = 8'h0f;
vram[12'h554] = 8'h0f;
vram[12'h555] = 8'h0f;
vram[12'h556] = 8'h0f;
vram[12'h557] = 8'h0f;
vram[12'h558] = 8'h0f;
vram[12'h559] = 8'h0f;
vram[12'h55a] = 8'h0f;
vram[12'h55b] = 8'h0f;
vram[12'h55c] = 8'h0f;
vram[12'h55d] = 8'h0f;
vram[12'h55e] = 8'h0f;
vram[12'h55f] = 8'h0f;
vram[12'h560] = 8'h0f;
vram[12'h561] = 8'h0f;
vram[12'h562] = 8'h0f;
vram[12'h563] = 8'h0f;
vram[12'h564] = 8'h0f;
vram[12'h565] = 8'h0f;
vram[12'h566] = 8'h0f;
vram[12'h567] = 8'h0f;
vram[12'h568] = 8'h0f;
vram[12'h569] = 8'h0f;
vram[12'h56a] = 8'h0f;
vram[12'h56b] = 8'h0f;
vram[12'h56c] = 8'h0f;
vram[12'h56d] = 8'h0f;
vram[12'h56e] = 8'h0f;
vram[12'h56f] = 8'h0f;
vram[12'h570] = 8'h0f;
vram[12'h571] = 8'h0f;
vram[12'h572] = 8'h0f;
vram[12'h573] = 8'h0f;
vram[12'h574] = 8'h0f;
vram[12'h575] = 8'h0f;
vram[12'h576] = 8'h0f;
vram[12'h577] = 8'h0f;
vram[12'h578] = 8'h0f;
vram[12'h579] = 8'h0f;
vram[12'h57a] = 8'h0f;
vram[12'h57b] = 8'h0f;
vram[12'h57c] = 8'h0f;
vram[12'h57d] = 8'h0f;
vram[12'h57e] = 8'h0f;
vram[12'h57f] = 8'h0f;
vram[12'h580] = 8'h0f;
vram[12'h581] = 8'h0f;
vram[12'h582] = 8'h0f;
vram[12'h583] = 8'h0f;
vram[12'h584] = 8'h0f;
vram[12'h585] = 8'h0f;
vram[12'h586] = 8'h0f;
vram[12'h587] = 8'h0f;
vram[12'h588] = 8'h0f;
vram[12'h589] = 8'h0f;
vram[12'h58a] = 8'h0f;
vram[12'h58b] = 8'h0f;
vram[12'h58c] = 8'h0f;
vram[12'h58d] = 8'h0f;
vram[12'h58e] = 8'h0f;
vram[12'h58f] = 8'h0f;
vram[12'h590] = 8'h0f;
vram[12'h591] = 8'h0f;
vram[12'h592] = 8'h0f;
vram[12'h593] = 8'h0f;
vram[12'h594] = 8'h0f;
vram[12'h595] = 8'h0f;
vram[12'h596] = 8'h0f;
vram[12'h597] = 8'h0f;
vram[12'h598] = 8'h0f;
vram[12'h599] = 8'h0f;
vram[12'h59a] = 8'h0f;
vram[12'h59b] = 8'h0f;
vram[12'h59c] = 8'h0f;
vram[12'h59d] = 8'h0f;
vram[12'h59e] = 8'h0f;
vram[12'h59f] = 8'h0f;
vram[12'h5a0] = 8'h0f;
vram[12'h5a1] = 8'h0f;
vram[12'h5a2] = 8'h0f;
vram[12'h5a3] = 8'h0f;
vram[12'h5a4] = 8'h0f;
vram[12'h5a5] = 8'h0f;
vram[12'h5a6] = 8'h0f;
vram[12'h5a7] = 8'h0f;
vram[12'h5a8] = 8'h0f;
vram[12'h5a9] = 8'h0f;
vram[12'h5aa] = 8'h0f;
vram[12'h5ab] = 8'h0f;
vram[12'h5ac] = 8'h0f;
vram[12'h5ad] = 8'h0f;
vram[12'h5ae] = 8'h0f;
vram[12'h5af] = 8'h0f;
vram[12'h5b0] = 8'h0f;
vram[12'h5b1] = 8'h0f;
vram[12'h5b2] = 8'h0f;
vram[12'h5b3] = 8'h0f;
vram[12'h5b4] = 8'h0f;
vram[12'h5b5] = 8'h0f;
vram[12'h5b6] = 8'h0f;
vram[12'h5b7] = 8'h0f;
vram[12'h5b8] = 8'h0f;
vram[12'h5b9] = 8'h0f;
vram[12'h5ba] = 8'h0f;
vram[12'h5bb] = 8'h0f;
vram[12'h5bc] = 8'h0f;
vram[12'h5bd] = 8'h0f;
vram[12'h5be] = 8'h0f;
vram[12'h5bf] = 8'h0f;
vram[12'h5c0] = 8'h0f;
vram[12'h5c1] = 8'h0f;
vram[12'h5c2] = 8'h0f;
vram[12'h5c3] = 8'h0f;
vram[12'h5c4] = 8'h0f;
vram[12'h5c5] = 8'h0f;
vram[12'h5c6] = 8'h0f;
vram[12'h5c7] = 8'h0f;
vram[12'h5c8] = 8'h0f;
vram[12'h5c9] = 8'h0f;
vram[12'h5ca] = 8'h0f;
vram[12'h5cb] = 8'h0f;
vram[12'h5cc] = 8'h0f;
vram[12'h5cd] = 8'h0f;
vram[12'h5ce] = 8'h0f;
vram[12'h5cf] = 8'h0f;
vram[12'h5d0] = 8'h0f;
vram[12'h5d1] = 8'h0f;
vram[12'h5d2] = 8'h0f;
vram[12'h5d3] = 8'h0f;
vram[12'h5d4] = 8'h0f;
vram[12'h5d5] = 8'h0f;
vram[12'h5d6] = 8'h0f;
vram[12'h5d7] = 8'h0f;
vram[12'h5d8] = 8'h0f;
vram[12'h5d9] = 8'h0f;
vram[12'h5da] = 8'h0f;
vram[12'h5db] = 8'h0f;
vram[12'h5dc] = 8'h0f;
vram[12'h5dd] = 8'h0f;
vram[12'h5de] = 8'h0f;
vram[12'h5df] = 8'h0f;
vram[12'h5e0] = 8'h0f;
vram[12'h5e1] = 8'h0f;
vram[12'h5e2] = 8'h0f;
vram[12'h5e3] = 8'h0f;
vram[12'h5e4] = 8'h0f;
vram[12'h5e5] = 8'h0f;
vram[12'h5e6] = 8'h0f;
vram[12'h5e7] = 8'h0f;
vram[12'h5e8] = 8'h0f;
vram[12'h5e9] = 8'h0f;
vram[12'h5ea] = 8'h0f;
vram[12'h5eb] = 8'h0f;
vram[12'h5ec] = 8'h0f;
vram[12'h5ed] = 8'h0f;
vram[12'h5ee] = 8'h0f;
vram[12'h5ef] = 8'h0f;
vram[12'h5f0] = 8'h0f;
vram[12'h5f1] = 8'h0f;
vram[12'h5f2] = 8'h0f;
vram[12'h5f3] = 8'h0f;
vram[12'h5f4] = 8'h0f;
vram[12'h5f5] = 8'h0f;
vram[12'h5f6] = 8'h0f;
vram[12'h5f7] = 8'h0f;
vram[12'h5f8] = 8'h0f;
vram[12'h5f9] = 8'h0f;
vram[12'h5fa] = 8'h0f;
vram[12'h5fb] = 8'h0f;
vram[12'h5fc] = 8'h0f;
vram[12'h5fd] = 8'h0f;
vram[12'h5fe] = 8'h0f;
vram[12'h5ff] = 8'h0f;
vram[12'h600] = 8'h0f;
vram[12'h601] = 8'h0f;
vram[12'h602] = 8'h0f;
vram[12'h603] = 8'h0f;
vram[12'h604] = 8'h0f;
vram[12'h605] = 8'h0f;
vram[12'h606] = 8'h0f;
vram[12'h607] = 8'h0f;
vram[12'h608] = 8'h0f;
vram[12'h609] = 8'h0f;
vram[12'h60a] = 8'h0f;
vram[12'h60b] = 8'h0f;
vram[12'h60c] = 8'h0f;
vram[12'h60d] = 8'h0f;
vram[12'h60e] = 8'h0f;
vram[12'h60f] = 8'h0f;
vram[12'h610] = 8'h0f;
vram[12'h611] = 8'h0f;
vram[12'h612] = 8'h0f;
vram[12'h613] = 8'h0f;
vram[12'h614] = 8'h0f;
vram[12'h615] = 8'h0f;
vram[12'h616] = 8'h0f;
vram[12'h617] = 8'h0f;
vram[12'h618] = 8'h0f;
vram[12'h619] = 8'h0f;
vram[12'h61a] = 8'h0f;
vram[12'h61b] = 8'h0f;
vram[12'h61c] = 8'h0f;
vram[12'h61d] = 8'h0f;
vram[12'h61e] = 8'h0f;
vram[12'h61f] = 8'h0f;
vram[12'h620] = 8'h0f;
vram[12'h621] = 8'h0f;
vram[12'h622] = 8'h0f;
vram[12'h623] = 8'h0f;
vram[12'h624] = 8'h0f;
vram[12'h625] = 8'h0f;
vram[12'h626] = 8'h0f;
vram[12'h627] = 8'h0f;
vram[12'h628] = 8'h0f;
vram[12'h629] = 8'h0f;
vram[12'h62a] = 8'h0f;
vram[12'h62b] = 8'h0f;
vram[12'h62c] = 8'h0f;
vram[12'h62d] = 8'h0f;
vram[12'h62e] = 8'h0f;
vram[12'h62f] = 8'h0f;
vram[12'h630] = 8'h0f;
vram[12'h631] = 8'h0f;
vram[12'h632] = 8'h0f;
vram[12'h633] = 8'h0f;
vram[12'h634] = 8'h0f;
vram[12'h635] = 8'h0f;
vram[12'h636] = 8'h0f;
vram[12'h637] = 8'h0f;
vram[12'h638] = 8'h0f;
vram[12'h639] = 8'h0f;
vram[12'h63a] = 8'h0f;
vram[12'h63b] = 8'h0f;
vram[12'h63c] = 8'h0f;
vram[12'h63d] = 8'h0f;
vram[12'h63e] = 8'h0f;
vram[12'h63f] = 8'h0f;
vram[12'h640] = 8'h0f;
vram[12'h641] = 8'h0f;
vram[12'h642] = 8'h0f;
vram[12'h643] = 8'h0f;
vram[12'h644] = 8'h0f;
vram[12'h645] = 8'h0f;
vram[12'h646] = 8'h0f;
vram[12'h647] = 8'h0f;
vram[12'h648] = 8'h0f;
vram[12'h649] = 8'h0f;
vram[12'h64a] = 8'h0f;
vram[12'h64b] = 8'h0f;
vram[12'h64c] = 8'h0f;
vram[12'h64d] = 8'h0f;
vram[12'h64e] = 8'h0f;
vram[12'h64f] = 8'h0f;
vram[12'h650] = 8'h0f;
vram[12'h651] = 8'h0f;
vram[12'h652] = 8'h0f;
vram[12'h653] = 8'h0f;
vram[12'h654] = 8'h0f;
vram[12'h655] = 8'h0f;
vram[12'h656] = 8'h0f;
vram[12'h657] = 8'h0f;
vram[12'h658] = 8'h0f;
vram[12'h659] = 8'h0f;
vram[12'h65a] = 8'h0f;
vram[12'h65b] = 8'h0f;
vram[12'h65c] = 8'h0f;
vram[12'h65d] = 8'h0f;
vram[12'h65e] = 8'h0f;
vram[12'h65f] = 8'h0f;
vram[12'h660] = 8'h0f;
vram[12'h661] = 8'h0f;
vram[12'h662] = 8'h0f;
vram[12'h663] = 8'h0f;
vram[12'h664] = 8'h0f;
vram[12'h665] = 8'h0f;
vram[12'h666] = 8'h0f;
vram[12'h667] = 8'h0f;
vram[12'h668] = 8'h0f;
vram[12'h669] = 8'h0f;
vram[12'h66a] = 8'h0f;
vram[12'h66b] = 8'h0f;
vram[12'h66c] = 8'h0f;
vram[12'h66d] = 8'h0f;
vram[12'h66e] = 8'h0f;
vram[12'h66f] = 8'h0f;
vram[12'h670] = 8'h0f;
vram[12'h671] = 8'h0f;
vram[12'h672] = 8'h0f;
vram[12'h673] = 8'h0f;
vram[12'h674] = 8'h0f;
vram[12'h675] = 8'h0f;
vram[12'h676] = 8'h0f;
vram[12'h677] = 8'h0f;
vram[12'h678] = 8'h0f;
vram[12'h679] = 8'h0f;
vram[12'h67a] = 8'h0f;
vram[12'h67b] = 8'h0f;
vram[12'h67c] = 8'h0f;
vram[12'h67d] = 8'h0f;
vram[12'h67e] = 8'h0f;
vram[12'h67f] = 8'h0f;
vram[12'h680] = 8'h0f;
vram[12'h681] = 8'h0f;
vram[12'h682] = 8'h0f;
vram[12'h683] = 8'h0f;
vram[12'h684] = 8'h0f;
vram[12'h685] = 8'h0f;
vram[12'h686] = 8'h0f;
vram[12'h687] = 8'h0f;
vram[12'h688] = 8'h0f;
vram[12'h689] = 8'h0f;
vram[12'h68a] = 8'h0f;
vram[12'h68b] = 8'h0f;
vram[12'h68c] = 8'h0f;
vram[12'h68d] = 8'h0f;
vram[12'h68e] = 8'h0f;
vram[12'h68f] = 8'h0f;
vram[12'h690] = 8'h0f;
vram[12'h691] = 8'h0f;
vram[12'h692] = 8'h0f;
vram[12'h693] = 8'h0f;
vram[12'h694] = 8'h0f;
vram[12'h695] = 8'h0f;
vram[12'h696] = 8'h0f;
vram[12'h697] = 8'h0f;
vram[12'h698] = 8'h0f;
vram[12'h699] = 8'h0f;
vram[12'h69a] = 8'h0f;
vram[12'h69b] = 8'h0f;
vram[12'h69c] = 8'h0f;
vram[12'h69d] = 8'h0f;
vram[12'h69e] = 8'h0f;
vram[12'h69f] = 8'h0f;
vram[12'h6a0] = 8'h0f;
vram[12'h6a1] = 8'h0f;
vram[12'h6a2] = 8'h0f;
vram[12'h6a3] = 8'h0f;
vram[12'h6a4] = 8'h0f;
vram[12'h6a5] = 8'h0f;
vram[12'h6a6] = 8'h0f;
vram[12'h6a7] = 8'h0f;
vram[12'h6a8] = 8'h0f;
vram[12'h6a9] = 8'h0f;
vram[12'h6aa] = 8'h0f;
vram[12'h6ab] = 8'h0f;
vram[12'h6ac] = 8'h0f;
vram[12'h6ad] = 8'h0f;
vram[12'h6ae] = 8'h0f;
vram[12'h6af] = 8'h0f;
vram[12'h6b0] = 8'h0f;
vram[12'h6b1] = 8'h0f;
vram[12'h6b2] = 8'h0f;
vram[12'h6b3] = 8'h0f;
vram[12'h6b4] = 8'h0f;
vram[12'h6b5] = 8'h0f;
vram[12'h6b6] = 8'h0f;
vram[12'h6b7] = 8'h0f;
vram[12'h6b8] = 8'h0f;
vram[12'h6b9] = 8'h0f;
vram[12'h6ba] = 8'h0f;
vram[12'h6bb] = 8'h0f;
vram[12'h6bc] = 8'h0f;
vram[12'h6bd] = 8'h0f;
vram[12'h6be] = 8'h0f;
vram[12'h6bf] = 8'h0f;
vram[12'h6c0] = 8'h0f;
vram[12'h6c1] = 8'h0f;
vram[12'h6c2] = 8'h0f;
vram[12'h6c3] = 8'h0f;
vram[12'h6c4] = 8'h0f;
vram[12'h6c5] = 8'h0f;
vram[12'h6c6] = 8'h0f;
vram[12'h6c7] = 8'h0f;
vram[12'h6c8] = 8'h0f;
vram[12'h6c9] = 8'h0f;
vram[12'h6ca] = 8'h0f;
vram[12'h6cb] = 8'h0f;
vram[12'h6cc] = 8'h0f;
vram[12'h6cd] = 8'h0f;
vram[12'h6ce] = 8'h0f;
vram[12'h6cf] = 8'h0f;
vram[12'h6d0] = 8'h0f;
vram[12'h6d1] = 8'h0f;
vram[12'h6d2] = 8'h0f;
vram[12'h6d3] = 8'h0f;
vram[12'h6d4] = 8'h0f;
vram[12'h6d5] = 8'h0f;
vram[12'h6d6] = 8'h0f;
vram[12'h6d7] = 8'h0f;
vram[12'h6d8] = 8'h0f;
vram[12'h6d9] = 8'h0f;
vram[12'h6da] = 8'h0f;
vram[12'h6db] = 8'h0f;
vram[12'h6dc] = 8'h0f;
vram[12'h6dd] = 8'h0f;
vram[12'h6de] = 8'h0f;
vram[12'h6df] = 8'h0f;
vram[12'h6e0] = 8'h0f;
vram[12'h6e1] = 8'h0f;
vram[12'h6e2] = 8'h0f;
vram[12'h6e3] = 8'h0f;
vram[12'h6e4] = 8'h0f;
vram[12'h6e5] = 8'h0f;
vram[12'h6e6] = 8'h0f;
vram[12'h6e7] = 8'h0f;
vram[12'h6e8] = 8'h0f;
vram[12'h6e9] = 8'h0f;
vram[12'h6ea] = 8'h0f;
vram[12'h6eb] = 8'h0f;
vram[12'h6ec] = 8'h0f;
vram[12'h6ed] = 8'h0f;
vram[12'h6ee] = 8'h0f;
vram[12'h6ef] = 8'h0f;
vram[12'h6f0] = 8'h0f;
vram[12'h6f1] = 8'h0f;
vram[12'h6f2] = 8'h0f;
vram[12'h6f3] = 8'h0f;
vram[12'h6f4] = 8'h0f;
vram[12'h6f5] = 8'h0f;
vram[12'h6f6] = 8'h0f;
vram[12'h6f7] = 8'h0f;
vram[12'h6f8] = 8'h0f;
vram[12'h6f9] = 8'h0f;
vram[12'h6fa] = 8'h0f;
vram[12'h6fb] = 8'h0f;
vram[12'h6fc] = 8'h0f;
vram[12'h6fd] = 8'h0f;
vram[12'h6fe] = 8'h0f;
vram[12'h6ff] = 8'h0f;
vram[12'h700] = 8'h0f;
vram[12'h701] = 8'h0f;
vram[12'h702] = 8'h0f;
vram[12'h703] = 8'h0f;
vram[12'h704] = 8'h0f;
vram[12'h705] = 8'h0f;
vram[12'h706] = 8'h0f;
vram[12'h707] = 8'h0f;
vram[12'h708] = 8'h0f;
vram[12'h709] = 8'h0f;
vram[12'h70a] = 8'h0f;
vram[12'h70b] = 8'h0f;
vram[12'h70c] = 8'h0f;
vram[12'h70d] = 8'h0f;
vram[12'h70e] = 8'h0f;
vram[12'h70f] = 8'h0f;
vram[12'h710] = 8'h0f;
vram[12'h711] = 8'h0f;
vram[12'h712] = 8'h0f;
vram[12'h713] = 8'h0f;
vram[12'h714] = 8'h0f;
vram[12'h715] = 8'h0f;
vram[12'h716] = 8'h0f;
vram[12'h717] = 8'h0f;
vram[12'h718] = 8'h0f;
vram[12'h719] = 8'h0f;
vram[12'h71a] = 8'h0f;
vram[12'h71b] = 8'h0f;
vram[12'h71c] = 8'h0f;
vram[12'h71d] = 8'h0f;
vram[12'h71e] = 8'h0f;
vram[12'h71f] = 8'h0f;
vram[12'h720] = 8'h0f;
vram[12'h721] = 8'h0f;
vram[12'h722] = 8'h0f;
vram[12'h723] = 8'h0f;
vram[12'h724] = 8'h0f;
vram[12'h725] = 8'h0f;
vram[12'h726] = 8'h0f;
vram[12'h727] = 8'h0f;
vram[12'h728] = 8'h0f;
vram[12'h729] = 8'h0f;
vram[12'h72a] = 8'h0f;
vram[12'h72b] = 8'h0f;
vram[12'h72c] = 8'h0f;
vram[12'h72d] = 8'h0f;
vram[12'h72e] = 8'h0f;
vram[12'h72f] = 8'h0f;
vram[12'h730] = 8'h0f;
vram[12'h731] = 8'h0f;
vram[12'h732] = 8'h0f;
vram[12'h733] = 8'h0f;
vram[12'h734] = 8'h0f;
vram[12'h735] = 8'h0f;
vram[12'h736] = 8'h0f;
vram[12'h737] = 8'h0f;
vram[12'h738] = 8'h0f;
vram[12'h739] = 8'h0f;
vram[12'h73a] = 8'h0f;
vram[12'h73b] = 8'h0f;
vram[12'h73c] = 8'h0f;
vram[12'h73d] = 8'h0f;
vram[12'h73e] = 8'h0f;
vram[12'h73f] = 8'h0f;
vram[12'h740] = 8'h0f;
vram[12'h741] = 8'h0f;
vram[12'h742] = 8'h0f;
vram[12'h743] = 8'h0f;
vram[12'h744] = 8'h0f;
vram[12'h745] = 8'h0f;
vram[12'h746] = 8'h0f;
vram[12'h747] = 8'h0f;
vram[12'h748] = 8'h0f;
vram[12'h749] = 8'h0f;
vram[12'h74a] = 8'h0f;
vram[12'h74b] = 8'h0f;
vram[12'h74c] = 8'h0f;
vram[12'h74d] = 8'h0f;
vram[12'h74e] = 8'h0f;
vram[12'h74f] = 8'h0f;
vram[12'h750] = 8'h0f;
vram[12'h751] = 8'h0f;
vram[12'h752] = 8'h0f;
vram[12'h753] = 8'h0f;
vram[12'h754] = 8'h0f;
vram[12'h755] = 8'h0f;
vram[12'h756] = 8'h0f;
vram[12'h757] = 8'h0f;
vram[12'h758] = 8'h0f;
vram[12'h759] = 8'h0f;
vram[12'h75a] = 8'h0f;
vram[12'h75b] = 8'h0f;
vram[12'h75c] = 8'h0f;
vram[12'h75d] = 8'h0f;
vram[12'h75e] = 8'h0f;
vram[12'h75f] = 8'h0f;
vram[12'h760] = 8'h0f;
vram[12'h761] = 8'h0f;
vram[12'h762] = 8'h0f;
vram[12'h763] = 8'h0f;
vram[12'h764] = 8'h0f;
vram[12'h765] = 8'h0f;
vram[12'h766] = 8'h0f;
vram[12'h767] = 8'h0f;
vram[12'h768] = 8'h0f;
vram[12'h769] = 8'h0f;
vram[12'h76a] = 8'h0f;
vram[12'h76b] = 8'h0f;
vram[12'h76c] = 8'h0f;
vram[12'h76d] = 8'h0f;
vram[12'h76e] = 8'h0f;
vram[12'h76f] = 8'h0f;
vram[12'h770] = 8'h0f;
vram[12'h771] = 8'h0f;
vram[12'h772] = 8'h0f;
vram[12'h773] = 8'h0f;
vram[12'h774] = 8'h0f;
vram[12'h775] = 8'h0f;
vram[12'h776] = 8'h0f;
vram[12'h777] = 8'h0f;
vram[12'h778] = 8'h0f;
vram[12'h779] = 8'h0f;
vram[12'h77a] = 8'h0f;
vram[12'h77b] = 8'h0f;
vram[12'h77c] = 8'h0f;
vram[12'h77d] = 8'h0f;
vram[12'h77e] = 8'h0f;
vram[12'h77f] = 8'h0f;
vram[12'h780] = 8'h0f;
vram[12'h781] = 8'h0f;
vram[12'h782] = 8'h0f;
vram[12'h783] = 8'h0f;
vram[12'h784] = 8'h0f;
vram[12'h785] = 8'h0f;
vram[12'h786] = 8'h0f;
vram[12'h787] = 8'h0f;
vram[12'h788] = 8'h0f;
vram[12'h789] = 8'h0f;
vram[12'h78a] = 8'h0f;
vram[12'h78b] = 8'h0f;
vram[12'h78c] = 8'h0f;
vram[12'h78d] = 8'h0f;
vram[12'h78e] = 8'h0f;
vram[12'h78f] = 8'h0f;
vram[12'h790] = 8'h0f;
vram[12'h791] = 8'h0f;
vram[12'h792] = 8'h0f;
vram[12'h793] = 8'h0f;
vram[12'h794] = 8'h0f;
vram[12'h795] = 8'h0f;
vram[12'h796] = 8'h0f;
vram[12'h797] = 8'h0f;
vram[12'h798] = 8'h0f;
vram[12'h799] = 8'h0f;
vram[12'h79a] = 8'h0f;
vram[12'h79b] = 8'h0f;
vram[12'h79c] = 8'h0f;
vram[12'h79d] = 8'h0f;
vram[12'h79e] = 8'h0f;
vram[12'h79f] = 8'h0f;
vram[12'h7a0] = 8'h0f;
vram[12'h7a1] = 8'h0f;
vram[12'h7a2] = 8'h0f;
vram[12'h7a3] = 8'h0f;
vram[12'h7a4] = 8'h0f;
vram[12'h7a5] = 8'h0f;
vram[12'h7a6] = 8'h0f;
vram[12'h7a7] = 8'h0f;
vram[12'h7a8] = 8'h0f;
vram[12'h7a9] = 8'h0f;
vram[12'h7aa] = 8'h0f;
vram[12'h7ab] = 8'h0f;
vram[12'h7ac] = 8'h0f;
vram[12'h7ad] = 8'h0f;
vram[12'h7ae] = 8'h0f;
vram[12'h7af] = 8'h0f;
vram[12'h7b0] = 8'h0f;
vram[12'h7b1] = 8'h0f;
vram[12'h7b2] = 8'h0f;
vram[12'h7b3] = 8'h0f;
vram[12'h7b4] = 8'h0f;
vram[12'h7b5] = 8'h0f;
vram[12'h7b6] = 8'h0f;
vram[12'h7b7] = 8'h0f;
vram[12'h7b8] = 8'h0f;
vram[12'h7b9] = 8'h0f;
vram[12'h7ba] = 8'h0f;
vram[12'h7bb] = 8'h0f;
vram[12'h7bc] = 8'h0f;
vram[12'h7bd] = 8'h0f;
vram[12'h7be] = 8'h0f;
vram[12'h7bf] = 8'h0f;
vram[12'h7c0] = 8'h0f;
vram[12'h7c1] = 8'h0f;
vram[12'h7c2] = 8'h0f;
vram[12'h7c3] = 8'h0f;
vram[12'h7c4] = 8'h0f;
vram[12'h7c5] = 8'h0f;
vram[12'h7c6] = 8'h0f;
vram[12'h7c7] = 8'h0f;
vram[12'h7c8] = 8'h0f;
vram[12'h7c9] = 8'h0f;
vram[12'h7ca] = 8'h0f;
vram[12'h7cb] = 8'h0f;
vram[12'h7cc] = 8'h0f;
vram[12'h7cd] = 8'h0f;
vram[12'h7ce] = 8'h0f;
vram[12'h7cf] = 8'h0f;
vram[12'h7d0] = 8'h0f;
vram[12'h7d1] = 8'h0f;
vram[12'h7d2] = 8'h0f;
vram[12'h7d3] = 8'h0f;
vram[12'h7d4] = 8'h0f;
vram[12'h7d5] = 8'h0f;
vram[12'h7d6] = 8'h0f;
vram[12'h7d7] = 8'h0f;
vram[12'h7d8] = 8'h0f;
vram[12'h7d9] = 8'h0f;
vram[12'h7da] = 8'h0f;
vram[12'h7db] = 8'h0f;
vram[12'h7dc] = 8'h0f;
vram[12'h7dd] = 8'h0f;
vram[12'h7de] = 8'h0f;
vram[12'h7df] = 8'h0f;
vram[12'h7e0] = 8'h0f;
vram[12'h7e1] = 8'h0f;
vram[12'h7e2] = 8'h0f;
vram[12'h7e3] = 8'h0f;
vram[12'h7e4] = 8'h0f;
vram[12'h7e5] = 8'h0f;
vram[12'h7e6] = 8'h0f;
vram[12'h7e7] = 8'h0f;
vram[12'h7e8] = 8'h0f;
vram[12'h7e9] = 8'h0f;
vram[12'h7ea] = 8'h0f;
vram[12'h7eb] = 8'h0f;
vram[12'h7ec] = 8'h0f;
vram[12'h7ed] = 8'h0f;
vram[12'h7ee] = 8'h0f;
vram[12'h7ef] = 8'h0f;
vram[12'h7f0] = 8'h0f;
vram[12'h7f1] = 8'h0f;
vram[12'h7f2] = 8'h0f;
vram[12'h7f3] = 8'h0f;
vram[12'h7f4] = 8'h0f;
vram[12'h7f5] = 8'h0f;
vram[12'h7f6] = 8'h0f;
vram[12'h7f7] = 8'h0f;
vram[12'h7f8] = 8'h0f;
vram[12'h7f9] = 8'h0f;
vram[12'h7fa] = 8'h0f;
vram[12'h7fb] = 8'h0f;
vram[12'h7fc] = 8'h0f;
vram[12'h7fd] = 8'h0f;
vram[12'h7fe] = 8'h0f;
vram[12'h7ff] = 8'h0f;
vram[12'h800] = 8'h00;
vram[12'h801] = 8'h00;
vram[12'h802] = 8'h00;
vram[12'h803] = 8'h00;
vram[12'h804] = 8'h00;
vram[12'h805] = 8'h00;
vram[12'h806] = 8'h00;
vram[12'h807] = 8'h00;
vram[12'h808] = 8'h01;
vram[12'h809] = 8'h03;
vram[12'h80a] = 8'h03;
vram[12'h80b] = 8'h06;
vram[12'h80c] = 8'h06;
vram[12'h80d] = 8'h0c;
vram[12'h80e] = 8'h0c;
vram[12'h80f] = 8'h18;
vram[12'h810] = 8'he0;
vram[12'h811] = 8'h38;
vram[12'h812] = 8'h0e;
vram[12'h813] = 8'h03;
vram[12'h814] = 8'h0e;
vram[12'h815] = 8'h38;
vram[12'h816] = 8'he0;
vram[12'h817] = 8'h00;
vram[12'h818] = 8'h07;
vram[12'h819] = 8'h1c;
vram[12'h81a] = 8'h70;
vram[12'h81b] = 8'hc0;
vram[12'h81c] = 8'h30;
vram[12'h81d] = 8'h1c;
vram[12'h81e] = 8'h07;
vram[12'h81f] = 8'h00;
vram[12'h820] = 8'hc3;
vram[12'h821] = 8'hc3;
vram[12'h822] = 8'h66;
vram[12'h823] = 8'h66;
vram[12'h824] = 8'h3c;
vram[12'h825] = 8'h3c;
vram[12'h826] = 8'h18;
vram[12'h827] = 8'h18;
vram[12'h828] = 8'h18;
vram[12'h829] = 8'h18;
vram[12'h82a] = 8'h3c;
vram[12'h82b] = 8'h3c;
vram[12'h82c] = 8'h66;
vram[12'h82d] = 8'h66;
vram[12'h82e] = 8'hc3;
vram[12'h82f] = 8'hc3;
vram[12'h830] = 8'h00;
vram[12'h831] = 8'h00;
vram[12'h832] = 8'h00;
vram[12'h833] = 8'h10;
vram[12'h834] = 8'h00;
vram[12'h835] = 8'h00;
vram[12'h836] = 8'h00;
vram[12'h837] = 8'h00;
vram[12'h838] = 8'h00;
vram[12'h839] = 8'h3f;
vram[12'h83a] = 8'h3f;
vram[12'h83b] = 8'h3f;
vram[12'h83c] = 8'h3f;
vram[12'h83d] = 8'h3f;
vram[12'h83e] = 8'h3f;
vram[12'h83f] = 8'h00;
vram[12'h840] = 8'h00;
vram[12'h841] = 8'hfc;
vram[12'h842] = 8'hfc;
vram[12'h843] = 8'hfc;
vram[12'h844] = 8'hfc;
vram[12'h845] = 8'hfc;
vram[12'h846] = 8'hfc;
vram[12'h847] = 8'h00;
vram[12'h848] = 8'h00;
vram[12'h849] = 8'h54;
vram[12'h84a] = 8'h2a;
vram[12'h84b] = 8'h54;
vram[12'h84c] = 8'h2a;
vram[12'h84d] = 8'h54;
vram[12'h84e] = 8'h2a;
vram[12'h84f] = 8'h00;
vram[12'h850] = 8'h00;
vram[12'h851] = 8'h00;
vram[12'h852] = 8'h18;
vram[12'h853] = 8'h3c;
vram[12'h854] = 8'h3c;
vram[12'h855] = 8'h7e;
vram[12'h856] = 8'h7e;
vram[12'h857] = 8'h7e;
vram[12'h858] = 8'h7e;
vram[12'h859] = 8'h7e;
vram[12'h85a] = 8'h7e;
vram[12'h85b] = 8'h3c;
vram[12'h85c] = 8'h3c;
vram[12'h85d] = 8'h18;
vram[12'h85e] = 8'h00;
vram[12'h85f] = 8'h00;
vram[12'h860] = 8'h07;
vram[12'h861] = 8'h1f;
vram[12'h862] = 8'h3f;
vram[12'h863] = 8'h7f;
vram[12'h864] = 8'h7f;
vram[12'h865] = 8'hff;
vram[12'h866] = 8'hff;
vram[12'h867] = 8'hff;
vram[12'h868] = 8'he0;
vram[12'h869] = 8'hf8;
vram[12'h86a] = 8'hfc;
vram[12'h86b] = 8'hfe;
vram[12'h86c] = 8'hfe;
vram[12'h86d] = 8'hff;
vram[12'h86e] = 8'hff;
vram[12'h86f] = 8'hff;
vram[12'h870] = 8'hff;
vram[12'h871] = 8'hff;
vram[12'h872] = 8'hff;
vram[12'h873] = 8'hfe;
vram[12'h874] = 8'hfe;
vram[12'h875] = 8'hfc;
vram[12'h876] = 8'hf8;
vram[12'h877] = 8'he0;
vram[12'h878] = 8'hff;
vram[12'h879] = 8'hff;
vram[12'h87a] = 8'hff;
vram[12'h87b] = 8'h7f;
vram[12'h87c] = 8'h7f;
vram[12'h87d] = 8'h3f;
vram[12'h87e] = 8'h1f;
vram[12'h87f] = 8'h07;
vram[12'h880] = 8'h24;
vram[12'h881] = 8'h42;
vram[12'h882] = 8'h81;
vram[12'h883] = 8'h00;
vram[12'h884] = 8'h00;
vram[12'h885] = 8'h81;
vram[12'h886] = 8'h42;
vram[12'h887] = 8'h24;
vram[12'h888] = 8'h00;
vram[12'h889] = 8'h00;
vram[12'h88a] = 8'h02;
vram[12'h88b] = 8'h00;
vram[12'h88c] = 8'h00;
vram[12'h88d] = 8'h00;
vram[12'h88e] = 8'h20;
vram[12'h88f] = 8'h00;
vram[12'h890] = 8'h20;
vram[12'h891] = 8'h00;
vram[12'h892] = 8'h02;
vram[12'h893] = 8'h00;
vram[12'h894] = 8'h20;
vram[12'h895] = 8'h00;
vram[12'h896] = 8'h02;
vram[12'h897] = 8'h00;
vram[12'h898] = 8'h22;
vram[12'h899] = 8'h00;
vram[12'h89a] = 8'h88;
vram[12'h89b] = 8'h00;
vram[12'h89c] = 8'h22;
vram[12'h89d] = 8'h00;
vram[12'h89e] = 8'h88;
vram[12'h89f] = 8'h00;
vram[12'h8a0] = 8'h88;
vram[12'h8a1] = 8'h00;
vram[12'h8a2] = 8'h55;
vram[12'h8a3] = 8'h00;
vram[12'h8a4] = 8'h22;
vram[12'h8a5] = 8'h00;
vram[12'h8a6] = 8'h55;
vram[12'h8a7] = 8'h00;
vram[12'h8a8] = 8'hff;
vram[12'h8a9] = 8'hbb;
vram[12'h8aa] = 8'hff;
vram[12'h8ab] = 8'hee;
vram[12'h8ac] = 8'hff;
vram[12'h8ad] = 8'hbb;
vram[12'h8ae] = 8'hff;
vram[12'h8af] = 8'hee;
vram[12'h8b0] = 8'hbf;
vram[12'h8b1] = 8'hff;
vram[12'h8b2] = 8'hfb;
vram[12'h8b3] = 8'hff;
vram[12'h8b4] = 8'hbf;
vram[12'h8b5] = 8'hff;
vram[12'h8b6] = 8'hfb;
vram[12'h8b7] = 8'hff;
vram[12'h8b8] = 8'hff;
vram[12'h8b9] = 8'hff;
vram[12'h8ba] = 8'hdf;
vram[12'h8bb] = 8'hff;
vram[12'h8bc] = 8'hff;
vram[12'h8bd] = 8'hff;
vram[12'h8be] = 8'hfd;
vram[12'h8bf] = 8'hff;
vram[12'h8c0] = 8'haa;
vram[12'h8c1] = 8'h00;
vram[12'h8c2] = 8'haa;
vram[12'h8c3] = 8'h00;
vram[12'h8c4] = 8'haa;
vram[12'h8c5] = 8'h00;
vram[12'h8c6] = 8'haa;
vram[12'h8c7] = 8'h00;
vram[12'h8c8] = 8'h00;
vram[12'h8c9] = 8'h44;
vram[12'h8ca] = 8'h00;
vram[12'h8cb] = 8'h00;
vram[12'h8cc] = 8'h00;
vram[12'h8cd] = 8'h44;
vram[12'h8ce] = 8'h00;
vram[12'h8cf] = 8'h00;
vram[12'h8d0] = 8'hcc;
vram[12'h8d1] = 8'hcc;
vram[12'h8d2] = 8'h33;
vram[12'h8d3] = 8'h33;
vram[12'h8d4] = 8'hcc;
vram[12'h8d5] = 8'hcc;
vram[12'h8d6] = 8'h33;
vram[12'h8d7] = 8'h33;
vram[12'h8d8] = 8'h3c;
vram[12'h8d9] = 8'h66;
vram[12'h8da] = 8'h66;
vram[12'h8db] = 8'h30;
vram[12'h8dc] = 8'h18;
vram[12'h8dd] = 8'h00;
vram[12'h8de] = 8'h18;
vram[12'h8df] = 8'h00;
vram[12'h8e0] = 8'h33;
vram[12'h8e1] = 8'h66;
vram[12'h8e2] = 8'hcc;
vram[12'h8e3] = 8'h99;
vram[12'h8e4] = 8'h33;
vram[12'h8e5] = 8'h66;
vram[12'h8e6] = 8'hcc;
vram[12'h8e7] = 8'h99;
vram[12'h8e8] = 8'hcc;
vram[12'h8e9] = 8'h66;
vram[12'h8ea] = 8'h33;
vram[12'h8eb] = 8'h99;
vram[12'h8ec] = 8'hcc;
vram[12'h8ed] = 8'h66;
vram[12'h8ee] = 8'h33;
vram[12'h8ef] = 8'h99;
vram[12'h8f0] = 8'he0;
vram[12'h8f1] = 8'ha0;
vram[12'h8f2] = 8'hee;
vram[12'h8f3] = 8'hc8;
vram[12'h8f4] = 8'hae;
vram[12'h8f5] = 8'h02;
vram[12'h8f6] = 8'h0e;
vram[12'h8f7] = 8'h00;
vram[12'h8f8] = 8'ha0;
vram[12'h8f9] = 8'ha0;
vram[12'h8fa] = 8'hae;
vram[12'h8fb] = 8'ha8;
vram[12'h8fc] = 8'hee;
vram[12'h8fd] = 8'h02;
vram[12'h8fe] = 8'h0e;
vram[12'h8ff] = 8'h00;
vram[12'h900] = 8'h00;
vram[12'h901] = 8'h00;
vram[12'h902] = 8'h00;
vram[12'h903] = 8'h00;
vram[12'h904] = 8'h00;
vram[12'h905] = 8'h00;
vram[12'h906] = 8'h00;
vram[12'h907] = 8'h00;
vram[12'h908] = 8'h18;
vram[12'h909] = 8'h18;
vram[12'h90a] = 8'h18;
vram[12'h90b] = 8'h18;
vram[12'h90c] = 8'h18;
vram[12'h90d] = 8'h00;
vram[12'h90e] = 8'h18;
vram[12'h90f] = 8'h00;
vram[12'h910] = 8'h66;
vram[12'h911] = 8'h66;
vram[12'h912] = 8'h66;
vram[12'h913] = 8'h00;
vram[12'h914] = 8'h00;
vram[12'h915] = 8'h00;
vram[12'h916] = 8'h00;
vram[12'h917] = 8'h00;
vram[12'h918] = 8'h6c;
vram[12'h919] = 8'h6c;
vram[12'h91a] = 8'hfe;
vram[12'h91b] = 8'h6c;
vram[12'h91c] = 8'hfe;
vram[12'h91d] = 8'h6c;
vram[12'h91e] = 8'h6c;
vram[12'h91f] = 8'h00;
vram[12'h920] = 8'h18;
vram[12'h921] = 8'h3e;
vram[12'h922] = 8'h60;
vram[12'h923] = 8'h3c;
vram[12'h924] = 8'h06;
vram[12'h925] = 8'h7c;
vram[12'h926] = 8'h18;
vram[12'h927] = 8'h00;
vram[12'h928] = 8'h00;
vram[12'h929] = 8'hc6;
vram[12'h92a] = 8'hcc;
vram[12'h92b] = 8'h18;
vram[12'h92c] = 8'h30;
vram[12'h92d] = 8'h66;
vram[12'h92e] = 8'hc6;
vram[12'h92f] = 8'h00;
vram[12'h930] = 8'h38;
vram[12'h931] = 8'h6c;
vram[12'h932] = 8'h38;
vram[12'h933] = 8'h76;
vram[12'h934] = 8'hdc;
vram[12'h935] = 8'hcc;
vram[12'h936] = 8'h76;
vram[12'h937] = 8'h00;
vram[12'h938] = 8'h18;
vram[12'h939] = 8'h18;
vram[12'h93a] = 8'h30;
vram[12'h93b] = 8'h00;
vram[12'h93c] = 8'h00;
vram[12'h93d] = 8'h00;
vram[12'h93e] = 8'h00;
vram[12'h93f] = 8'h00;
vram[12'h940] = 8'h0c;
vram[12'h941] = 8'h18;
vram[12'h942] = 8'h30;
vram[12'h943] = 8'h30;
vram[12'h944] = 8'h30;
vram[12'h945] = 8'h18;
vram[12'h946] = 8'h0c;
vram[12'h947] = 8'h00;
vram[12'h948] = 8'h30;
vram[12'h949] = 8'h18;
vram[12'h94a] = 8'h0c;
vram[12'h94b] = 8'h0c;
vram[12'h94c] = 8'h0c;
vram[12'h94d] = 8'h18;
vram[12'h94e] = 8'h30;
vram[12'h94f] = 8'h00;
vram[12'h950] = 8'h00;
vram[12'h951] = 8'h66;
vram[12'h952] = 8'h3c;
vram[12'h953] = 8'hff;
vram[12'h954] = 8'h3c;
vram[12'h955] = 8'h66;
vram[12'h956] = 8'h00;
vram[12'h957] = 8'h00;
vram[12'h958] = 8'h00;
vram[12'h959] = 8'h18;
vram[12'h95a] = 8'h18;
vram[12'h95b] = 8'h7e;
vram[12'h95c] = 8'h18;
vram[12'h95d] = 8'h18;
vram[12'h95e] = 8'h00;
vram[12'h95f] = 8'h00;
vram[12'h960] = 8'h00;
vram[12'h961] = 8'h00;
vram[12'h962] = 8'h00;
vram[12'h963] = 8'h00;
vram[12'h964] = 8'h00;
vram[12'h965] = 8'h18;
vram[12'h966] = 8'h18;
vram[12'h967] = 8'h30;
vram[12'h968] = 8'h00;
vram[12'h969] = 8'h00;
vram[12'h96a] = 8'h00;
vram[12'h96b] = 8'h7e;
vram[12'h96c] = 8'h00;
vram[12'h96d] = 8'h00;
vram[12'h96e] = 8'h00;
vram[12'h96f] = 8'h00;
vram[12'h970] = 8'h00;
vram[12'h971] = 8'h00;
vram[12'h972] = 8'h00;
vram[12'h973] = 8'h00;
vram[12'h974] = 8'h00;
vram[12'h975] = 8'h18;
vram[12'h976] = 8'h18;
vram[12'h977] = 8'h00;
vram[12'h978] = 8'h03;
vram[12'h979] = 8'h06;
vram[12'h97a] = 8'h0c;
vram[12'h97b] = 8'h18;
vram[12'h97c] = 8'h30;
vram[12'h97d] = 8'h60;
vram[12'h97e] = 8'hc0;
vram[12'h97f] = 8'h00;
vram[12'h980] = 8'h3c;
vram[12'h981] = 8'h66;
vram[12'h982] = 8'h6e;
vram[12'h983] = 8'h76;
vram[12'h984] = 8'h66;
vram[12'h985] = 8'h66;
vram[12'h986] = 8'h3c;
vram[12'h987] = 8'h00;
vram[12'h988] = 8'h18;
vram[12'h989] = 8'h38;
vram[12'h98a] = 8'h18;
vram[12'h98b] = 8'h18;
vram[12'h98c] = 8'h18;
vram[12'h98d] = 8'h18;
vram[12'h98e] = 8'h7e;
vram[12'h98f] = 8'h00;
vram[12'h990] = 8'h3c;
vram[12'h991] = 8'h66;
vram[12'h992] = 8'h0c;
vram[12'h993] = 8'h18;
vram[12'h994] = 8'h30;
vram[12'h995] = 8'h60;
vram[12'h996] = 8'h7e;
vram[12'h997] = 8'h00;
vram[12'h998] = 8'h3c;
vram[12'h999] = 8'h66;
vram[12'h99a] = 8'h06;
vram[12'h99b] = 8'h1c;
vram[12'h99c] = 8'h06;
vram[12'h99d] = 8'h66;
vram[12'h99e] = 8'h3c;
vram[12'h99f] = 8'h00;
vram[12'h9a0] = 8'h1c;
vram[12'h9a1] = 8'h3c;
vram[12'h9a2] = 8'h6c;
vram[12'h9a3] = 8'hcc;
vram[12'h9a4] = 8'hfe;
vram[12'h9a5] = 8'h0c;
vram[12'h9a6] = 8'h0c;
vram[12'h9a7] = 8'h00;
vram[12'h9a8] = 8'h7e;
vram[12'h9a9] = 8'h60;
vram[12'h9aa] = 8'h7c;
vram[12'h9ab] = 8'h06;
vram[12'h9ac] = 8'h06;
vram[12'h9ad] = 8'h66;
vram[12'h9ae] = 8'h3c;
vram[12'h9af] = 8'h00;
vram[12'h9b0] = 8'h1c;
vram[12'h9b1] = 8'h30;
vram[12'h9b2] = 8'h60;
vram[12'h9b3] = 8'h7c;
vram[12'h9b4] = 8'h66;
vram[12'h9b5] = 8'h66;
vram[12'h9b6] = 8'h3c;
vram[12'h9b7] = 8'h00;
vram[12'h9b8] = 8'h7e;
vram[12'h9b9] = 8'h06;
vram[12'h9ba] = 8'h06;
vram[12'h9bb] = 8'h0c;
vram[12'h9bc] = 8'h18;
vram[12'h9bd] = 8'h18;
vram[12'h9be] = 8'h18;
vram[12'h9bf] = 8'h00;
vram[12'h9c0] = 8'h3c;
vram[12'h9c1] = 8'h66;
vram[12'h9c2] = 8'h66;
vram[12'h9c3] = 8'h3c;
vram[12'h9c4] = 8'h66;
vram[12'h9c5] = 8'h66;
vram[12'h9c6] = 8'h3c;
vram[12'h9c7] = 8'h00;
vram[12'h9c8] = 8'h3c;
vram[12'h9c9] = 8'h66;
vram[12'h9ca] = 8'h66;
vram[12'h9cb] = 8'h3e;
vram[12'h9cc] = 8'h06;
vram[12'h9cd] = 8'h0c;
vram[12'h9ce] = 8'h38;
vram[12'h9cf] = 8'h00;
vram[12'h9d0] = 8'h00;
vram[12'h9d1] = 8'h18;
vram[12'h9d2] = 8'h18;
vram[12'h9d3] = 8'h00;
vram[12'h9d4] = 8'h00;
vram[12'h9d5] = 8'h18;
vram[12'h9d6] = 8'h18;
vram[12'h9d7] = 8'h00;
vram[12'h9d8] = 8'h00;
vram[12'h9d9] = 8'h18;
vram[12'h9da] = 8'h18;
vram[12'h9db] = 8'h00;
vram[12'h9dc] = 8'h00;
vram[12'h9dd] = 8'h18;
vram[12'h9de] = 8'h18;
vram[12'h9df] = 8'h30;
vram[12'h9e0] = 8'h0c;
vram[12'h9e1] = 8'h18;
vram[12'h9e2] = 8'h30;
vram[12'h9e3] = 8'h60;
vram[12'h9e4] = 8'h30;
vram[12'h9e5] = 8'h18;
vram[12'h9e6] = 8'h0c;
vram[12'h9e7] = 8'h00;
vram[12'h9e8] = 8'h00;
vram[12'h9e9] = 8'h00;
vram[12'h9ea] = 8'h7e;
vram[12'h9eb] = 8'h00;
vram[12'h9ec] = 8'h7e;
vram[12'h9ed] = 8'h00;
vram[12'h9ee] = 8'h00;
vram[12'h9ef] = 8'h00;
vram[12'h9f0] = 8'h60;
vram[12'h9f1] = 8'h30;
vram[12'h9f2] = 8'h18;
vram[12'h9f3] = 8'h0c;
vram[12'h9f4] = 8'h18;
vram[12'h9f5] = 8'h30;
vram[12'h9f6] = 8'h60;
vram[12'h9f7] = 8'h00;
vram[12'h9f8] = 8'h3c;
vram[12'h9f9] = 8'h66;
vram[12'h9fa] = 8'h06;
vram[12'h9fb] = 8'h0c;
vram[12'h9fc] = 8'h18;
vram[12'h9fd] = 8'h00;
vram[12'h9fe] = 8'h18;
vram[12'h9ff] = 8'h00;
vram[12'ha00] = 8'h7c;
vram[12'ha01] = 8'hc6;
vram[12'ha02] = 8'hde;
vram[12'ha03] = 8'hde;
vram[12'ha04] = 8'hde;
vram[12'ha05] = 8'hc0;
vram[12'ha06] = 8'h7c;
vram[12'ha07] = 8'h00;
vram[12'ha08] = 8'h18;
vram[12'ha09] = 8'h3c;
vram[12'ha0a] = 8'h66;
vram[12'ha0b] = 8'h66;
vram[12'ha0c] = 8'h7e;
vram[12'ha0d] = 8'h66;
vram[12'ha0e] = 8'h66;
vram[12'ha0f] = 8'h00;
vram[12'ha10] = 8'h7c;
vram[12'ha11] = 8'h66;
vram[12'ha12] = 8'h66;
vram[12'ha13] = 8'h7c;
vram[12'ha14] = 8'h66;
vram[12'ha15] = 8'h66;
vram[12'ha16] = 8'h7c;
vram[12'ha17] = 8'h00;
vram[12'ha18] = 8'h3c;
vram[12'ha19] = 8'h66;
vram[12'ha1a] = 8'h60;
vram[12'ha1b] = 8'h60;
vram[12'ha1c] = 8'h60;
vram[12'ha1d] = 8'h66;
vram[12'ha1e] = 8'h3c;
vram[12'ha1f] = 8'h00;
vram[12'ha20] = 8'h78;
vram[12'ha21] = 8'h6c;
vram[12'ha22] = 8'h66;
vram[12'ha23] = 8'h66;
vram[12'ha24] = 8'h66;
vram[12'ha25] = 8'h6c;
vram[12'ha26] = 8'h78;
vram[12'ha27] = 8'h00;
vram[12'ha28] = 8'h7e;
vram[12'ha29] = 8'h60;
vram[12'ha2a] = 8'h60;
vram[12'ha2b] = 8'h7c;
vram[12'ha2c] = 8'h60;
vram[12'ha2d] = 8'h60;
vram[12'ha2e] = 8'h7e;
vram[12'ha2f] = 8'h00;
vram[12'ha30] = 8'h7e;
vram[12'ha31] = 8'h60;
vram[12'ha32] = 8'h60;
vram[12'ha33] = 8'h7c;
vram[12'ha34] = 8'h60;
vram[12'ha35] = 8'h60;
vram[12'ha36] = 8'h60;
vram[12'ha37] = 8'h00;
vram[12'ha38] = 8'h3c;
vram[12'ha39] = 8'h66;
vram[12'ha3a] = 8'h60;
vram[12'ha3b] = 8'h6e;
vram[12'ha3c] = 8'h66;
vram[12'ha3d] = 8'h66;
vram[12'ha3e] = 8'h3e;
vram[12'ha3f] = 8'h00;
vram[12'ha40] = 8'h66;
vram[12'ha41] = 8'h66;
vram[12'ha42] = 8'h66;
vram[12'ha43] = 8'h7e;
vram[12'ha44] = 8'h66;
vram[12'ha45] = 8'h66;
vram[12'ha46] = 8'h66;
vram[12'ha47] = 8'h00;
vram[12'ha48] = 8'h7e;
vram[12'ha49] = 8'h18;
vram[12'ha4a] = 8'h18;
vram[12'ha4b] = 8'h18;
vram[12'ha4c] = 8'h18;
vram[12'ha4d] = 8'h18;
vram[12'ha4e] = 8'h7e;
vram[12'ha4f] = 8'h00;
vram[12'ha50] = 8'h06;
vram[12'ha51] = 8'h06;
vram[12'ha52] = 8'h06;
vram[12'ha53] = 8'h06;
vram[12'ha54] = 8'h06;
vram[12'ha55] = 8'h66;
vram[12'ha56] = 8'h3c;
vram[12'ha57] = 8'h00;
vram[12'ha58] = 8'hc6;
vram[12'ha59] = 8'hcc;
vram[12'ha5a] = 8'hd8;
vram[12'ha5b] = 8'hf0;
vram[12'ha5c] = 8'hd8;
vram[12'ha5d] = 8'hcc;
vram[12'ha5e] = 8'hc6;
vram[12'ha5f] = 8'h00;
vram[12'ha60] = 8'h60;
vram[12'ha61] = 8'h60;
vram[12'ha62] = 8'h60;
vram[12'ha63] = 8'h60;
vram[12'ha64] = 8'h60;
vram[12'ha65] = 8'h60;
vram[12'ha66] = 8'h7e;
vram[12'ha67] = 8'h00;
vram[12'ha68] = 8'hc6;
vram[12'ha69] = 8'hee;
vram[12'ha6a] = 8'hfe;
vram[12'ha6b] = 8'hd6;
vram[12'ha6c] = 8'hc6;
vram[12'ha6d] = 8'hc6;
vram[12'ha6e] = 8'hc6;
vram[12'ha6f] = 8'h00;
vram[12'ha70] = 8'hc6;
vram[12'ha71] = 8'he6;
vram[12'ha72] = 8'hf6;
vram[12'ha73] = 8'hde;
vram[12'ha74] = 8'hce;
vram[12'ha75] = 8'hc6;
vram[12'ha76] = 8'hc6;
vram[12'ha77] = 8'h00;
vram[12'ha78] = 8'h3c;
vram[12'ha79] = 8'h66;
vram[12'ha7a] = 8'h66;
vram[12'ha7b] = 8'h66;
vram[12'ha7c] = 8'h66;
vram[12'ha7d] = 8'h66;
vram[12'ha7e] = 8'h3c;
vram[12'ha7f] = 8'h00;
vram[12'ha80] = 8'h7c;
vram[12'ha81] = 8'h66;
vram[12'ha82] = 8'h66;
vram[12'ha83] = 8'h7c;
vram[12'ha84] = 8'h60;
vram[12'ha85] = 8'h60;
vram[12'ha86] = 8'h60;
vram[12'ha87] = 8'h00;
vram[12'ha88] = 8'h3c;
vram[12'ha89] = 8'h66;
vram[12'ha8a] = 8'h66;
vram[12'ha8b] = 8'h66;
vram[12'ha8c] = 8'h66;
vram[12'ha8d] = 8'h6c;
vram[12'ha8e] = 8'h36;
vram[12'ha8f] = 8'h00;
vram[12'ha90] = 8'h7c;
vram[12'ha91] = 8'h66;
vram[12'ha92] = 8'h66;
vram[12'ha93] = 8'h7c;
vram[12'ha94] = 8'h6c;
vram[12'ha95] = 8'h66;
vram[12'ha96] = 8'h66;
vram[12'ha97] = 8'h00;
vram[12'ha98] = 8'h3c;
vram[12'ha99] = 8'h66;
vram[12'ha9a] = 8'h60;
vram[12'ha9b] = 8'h3c;
vram[12'ha9c] = 8'h06;
vram[12'ha9d] = 8'h66;
vram[12'ha9e] = 8'h3c;
vram[12'ha9f] = 8'h00;
vram[12'haa0] = 8'h7e;
vram[12'haa1] = 8'h18;
vram[12'haa2] = 8'h18;
vram[12'haa3] = 8'h18;
vram[12'haa4] = 8'h18;
vram[12'haa5] = 8'h18;
vram[12'haa6] = 8'h18;
vram[12'haa7] = 8'h00;
vram[12'haa8] = 8'h66;
vram[12'haa9] = 8'h66;
vram[12'haaa] = 8'h66;
vram[12'haab] = 8'h66;
vram[12'haac] = 8'h66;
vram[12'haad] = 8'h66;
vram[12'haae] = 8'h3c;
vram[12'haaf] = 8'h00;
vram[12'hab0] = 8'h66;
vram[12'hab1] = 8'h66;
vram[12'hab2] = 8'h66;
vram[12'hab3] = 8'h66;
vram[12'hab4] = 8'h66;
vram[12'hab5] = 8'h3c;
vram[12'hab6] = 8'h18;
vram[12'hab7] = 8'h00;
vram[12'hab8] = 8'hc6;
vram[12'hab9] = 8'hc6;
vram[12'haba] = 8'hc6;
vram[12'habb] = 8'hd6;
vram[12'habc] = 8'hfe;
vram[12'habd] = 8'hee;
vram[12'habe] = 8'hc6;
vram[12'habf] = 8'h00;
vram[12'hac0] = 8'hc3;
vram[12'hac1] = 8'h66;
vram[12'hac2] = 8'h3c;
vram[12'hac3] = 8'h18;
vram[12'hac4] = 8'h3c;
vram[12'hac5] = 8'h66;
vram[12'hac6] = 8'hc3;
vram[12'hac7] = 8'h00;
vram[12'hac8] = 8'hc3;
vram[12'hac9] = 8'h66;
vram[12'haca] = 8'h3c;
vram[12'hacb] = 8'h18;
vram[12'hacc] = 8'h18;
vram[12'hacd] = 8'h18;
vram[12'hace] = 8'h18;
vram[12'hacf] = 8'h00;
vram[12'had0] = 8'h7e;
vram[12'had1] = 8'h06;
vram[12'had2] = 8'h0c;
vram[12'had3] = 8'h18;
vram[12'had4] = 8'h30;
vram[12'had5] = 8'h60;
vram[12'had6] = 8'h7e;
vram[12'had7] = 8'h00;
vram[12'had8] = 8'h3c;
vram[12'had9] = 8'h30;
vram[12'hada] = 8'h30;
vram[12'hadb] = 8'h30;
vram[12'hadc] = 8'h30;
vram[12'hadd] = 8'h30;
vram[12'hade] = 8'h3c;
vram[12'hadf] = 8'h00;
vram[12'hae0] = 8'hc0;
vram[12'hae1] = 8'h60;
vram[12'hae2] = 8'h30;
vram[12'hae3] = 8'h18;
vram[12'hae4] = 8'h0c;
vram[12'hae5] = 8'h06;
vram[12'hae6] = 8'h03;
vram[12'hae7] = 8'h00;
vram[12'hae8] = 8'h3c;
vram[12'hae9] = 8'h0c;
vram[12'haea] = 8'h0c;
vram[12'haeb] = 8'h0c;
vram[12'haec] = 8'h0c;
vram[12'haed] = 8'h0c;
vram[12'haee] = 8'h3c;
vram[12'haef] = 8'h00;
vram[12'haf0] = 8'h10;
vram[12'haf1] = 8'h38;
vram[12'haf2] = 8'h6c;
vram[12'haf3] = 8'hc6;
vram[12'haf4] = 8'h00;
vram[12'haf5] = 8'h00;
vram[12'haf6] = 8'h00;
vram[12'haf7] = 8'h00;
vram[12'haf8] = 8'h00;
vram[12'haf9] = 8'h00;
vram[12'hafa] = 8'h00;
vram[12'hafb] = 8'h00;
vram[12'hafc] = 8'h00;
vram[12'hafd] = 8'h00;
vram[12'hafe] = 8'h00;
vram[12'haff] = 8'hff;
vram[12'hb00] = 8'h18;
vram[12'hb01] = 8'h0c;
vram[12'hb02] = 8'h06;
vram[12'hb03] = 8'h00;
vram[12'hb04] = 8'h00;
vram[12'hb05] = 8'h00;
vram[12'hb06] = 8'h00;
vram[12'hb07] = 8'h00;
vram[12'hb08] = 8'h00;
vram[12'hb09] = 8'h00;
vram[12'hb0a] = 8'h3c;
vram[12'hb0b] = 8'h06;
vram[12'hb0c] = 8'h3e;
vram[12'hb0d] = 8'h66;
vram[12'hb0e] = 8'h3e;
vram[12'hb0f] = 8'h00;
vram[12'hb10] = 8'h60;
vram[12'hb11] = 8'h60;
vram[12'hb12] = 8'h7c;
vram[12'hb13] = 8'h66;
vram[12'hb14] = 8'h66;
vram[12'hb15] = 8'h66;
vram[12'hb16] = 8'h7c;
vram[12'hb17] = 8'h00;
vram[12'hb18] = 8'h00;
vram[12'hb19] = 8'h00;
vram[12'hb1a] = 8'h3c;
vram[12'hb1b] = 8'h60;
vram[12'hb1c] = 8'h60;
vram[12'hb1d] = 8'h60;
vram[12'hb1e] = 8'h3c;
vram[12'hb1f] = 8'h00;
vram[12'hb20] = 8'h06;
vram[12'hb21] = 8'h06;
vram[12'hb22] = 8'h3e;
vram[12'hb23] = 8'h66;
vram[12'hb24] = 8'h66;
vram[12'hb25] = 8'h66;
vram[12'hb26] = 8'h3e;
vram[12'hb27] = 8'h00;
vram[12'hb28] = 8'h00;
vram[12'hb29] = 8'h00;
vram[12'hb2a] = 8'h3c;
vram[12'hb2b] = 8'h66;
vram[12'hb2c] = 8'h7e;
vram[12'hb2d] = 8'h60;
vram[12'hb2e] = 8'h3c;
vram[12'hb2f] = 8'h00;
vram[12'hb30] = 8'h1c;
vram[12'hb31] = 8'h30;
vram[12'hb32] = 8'h7c;
vram[12'hb33] = 8'h30;
vram[12'hb34] = 8'h30;
vram[12'hb35] = 8'h30;
vram[12'hb36] = 8'h30;
vram[12'hb37] = 8'h00;
vram[12'hb38] = 8'h00;
vram[12'hb39] = 8'h00;
vram[12'hb3a] = 8'h3e;
vram[12'hb3b] = 8'h66;
vram[12'hb3c] = 8'h66;
vram[12'hb3d] = 8'h3e;
vram[12'hb3e] = 8'h06;
vram[12'hb3f] = 8'h7c;
vram[12'hb40] = 8'h60;
vram[12'hb41] = 8'h60;
vram[12'hb42] = 8'h7c;
vram[12'hb43] = 8'h66;
vram[12'hb44] = 8'h66;
vram[12'hb45] = 8'h66;
vram[12'hb46] = 8'h66;
vram[12'hb47] = 8'h00;
vram[12'hb48] = 8'h18;
vram[12'hb49] = 8'h00;
vram[12'hb4a] = 8'h38;
vram[12'hb4b] = 8'h18;
vram[12'hb4c] = 8'h18;
vram[12'hb4d] = 8'h18;
vram[12'hb4e] = 8'h1e;
vram[12'hb4f] = 8'h00;
vram[12'hb50] = 8'h0c;
vram[12'hb51] = 8'h00;
vram[12'hb52] = 8'h0c;
vram[12'hb53] = 8'h0c;
vram[12'hb54] = 8'h0c;
vram[12'hb55] = 8'h0c;
vram[12'hb56] = 8'h0c;
vram[12'hb57] = 8'h78;
vram[12'hb58] = 8'h60;
vram[12'hb59] = 8'h60;
vram[12'hb5a] = 8'h66;
vram[12'hb5b] = 8'h6c;
vram[12'hb5c] = 8'h78;
vram[12'hb5d] = 8'h6c;
vram[12'hb5e] = 8'h66;
vram[12'hb5f] = 8'h00;
vram[12'hb60] = 8'h38;
vram[12'hb61] = 8'h18;
vram[12'hb62] = 8'h18;
vram[12'hb63] = 8'h18;
vram[12'hb64] = 8'h18;
vram[12'hb65] = 8'h18;
vram[12'hb66] = 8'h1e;
vram[12'hb67] = 8'h00;
vram[12'hb68] = 8'h00;
vram[12'hb69] = 8'h00;
vram[12'hb6a] = 8'hcc;
vram[12'hb6b] = 8'hfe;
vram[12'hb6c] = 8'hd6;
vram[12'hb6d] = 8'hd6;
vram[12'hb6e] = 8'hc6;
vram[12'hb6f] = 8'h00;
vram[12'hb70] = 8'h00;
vram[12'hb71] = 8'h00;
vram[12'hb72] = 8'h7c;
vram[12'hb73] = 8'h66;
vram[12'hb74] = 8'h66;
vram[12'hb75] = 8'h66;
vram[12'hb76] = 8'h66;
vram[12'hb77] = 8'h00;
vram[12'hb78] = 8'h00;
vram[12'hb79] = 8'h00;
vram[12'hb7a] = 8'h3c;
vram[12'hb7b] = 8'h66;
vram[12'hb7c] = 8'h66;
vram[12'hb7d] = 8'h66;
vram[12'hb7e] = 8'h3c;
vram[12'hb7f] = 8'h00;
vram[12'hb80] = 8'h00;
vram[12'hb81] = 8'h00;
vram[12'hb82] = 8'h7c;
vram[12'hb83] = 8'h66;
vram[12'hb84] = 8'h66;
vram[12'hb85] = 8'h7c;
vram[12'hb86] = 8'h60;
vram[12'hb87] = 8'h60;
vram[12'hb88] = 8'h00;
vram[12'hb89] = 8'h00;
vram[12'hb8a] = 8'h3e;
vram[12'hb8b] = 8'h66;
vram[12'hb8c] = 8'h66;
vram[12'hb8d] = 8'h3e;
vram[12'hb8e] = 8'h06;
vram[12'hb8f] = 8'h06;
vram[12'hb90] = 8'h00;
vram[12'hb91] = 8'h00;
vram[12'hb92] = 8'h7c;
vram[12'hb93] = 8'h66;
vram[12'hb94] = 8'h60;
vram[12'hb95] = 8'h60;
vram[12'hb96] = 8'h60;
vram[12'hb97] = 8'h00;
vram[12'hb98] = 8'h00;
vram[12'hb99] = 8'h00;
vram[12'hb9a] = 8'h3e;
vram[12'hb9b] = 8'h60;
vram[12'hb9c] = 8'h3c;
vram[12'hb9d] = 8'h06;
vram[12'hb9e] = 8'h7c;
vram[12'hb9f] = 8'h00;
vram[12'hba0] = 8'h30;
vram[12'hba1] = 8'h30;
vram[12'hba2] = 8'h7e;
vram[12'hba3] = 8'h30;
vram[12'hba4] = 8'h30;
vram[12'hba5] = 8'h30;
vram[12'hba6] = 8'h1e;
vram[12'hba7] = 8'h00;
vram[12'hba8] = 8'h00;
vram[12'hba9] = 8'h00;
vram[12'hbaa] = 8'h66;
vram[12'hbab] = 8'h66;
vram[12'hbac] = 8'h66;
vram[12'hbad] = 8'h66;
vram[12'hbae] = 8'h3e;
vram[12'hbaf] = 8'h00;
vram[12'hbb0] = 8'h00;
vram[12'hbb1] = 8'h00;
vram[12'hbb2] = 8'h66;
vram[12'hbb3] = 8'h66;
vram[12'hbb4] = 8'h66;
vram[12'hbb5] = 8'h3c;
vram[12'hbb6] = 8'h18;
vram[12'hbb7] = 8'h00;
vram[12'hbb8] = 8'h00;
vram[12'hbb9] = 8'h00;
vram[12'hbba] = 8'hc6;
vram[12'hbbb] = 8'hc6;
vram[12'hbbc] = 8'hd6;
vram[12'hbbd] = 8'h7c;
vram[12'hbbe] = 8'h6c;
vram[12'hbbf] = 8'h00;
vram[12'hbc0] = 8'h00;
vram[12'hbc1] = 8'h00;
vram[12'hbc2] = 8'hc6;
vram[12'hbc3] = 8'h6c;
vram[12'hbc4] = 8'h38;
vram[12'hbc5] = 8'h6c;
vram[12'hbc6] = 8'hc6;
vram[12'hbc7] = 8'h00;
vram[12'hbc8] = 8'h00;
vram[12'hbc9] = 8'h00;
vram[12'hbca] = 8'h66;
vram[12'hbcb] = 8'h66;
vram[12'hbcc] = 8'h66;
vram[12'hbcd] = 8'h3e;
vram[12'hbce] = 8'h06;
vram[12'hbcf] = 8'h3c;
vram[12'hbd0] = 8'h00;
vram[12'hbd1] = 8'h00;
vram[12'hbd2] = 8'h7e;
vram[12'hbd3] = 8'h0c;
vram[12'hbd4] = 8'h18;
vram[12'hbd5] = 8'h30;
vram[12'hbd6] = 8'h7e;
vram[12'hbd7] = 8'h00;
vram[12'hbd8] = 8'h0e;
vram[12'hbd9] = 8'h18;
vram[12'hbda] = 8'h18;
vram[12'hbdb] = 8'h70;
vram[12'hbdc] = 8'h18;
vram[12'hbdd] = 8'h18;
vram[12'hbde] = 8'h0e;
vram[12'hbdf] = 8'h00;
vram[12'hbe0] = 8'h18;
vram[12'hbe1] = 8'h18;
vram[12'hbe2] = 8'h18;
vram[12'hbe3] = 8'h18;
vram[12'hbe4] = 8'h18;
vram[12'hbe5] = 8'h18;
vram[12'hbe6] = 8'h18;
vram[12'hbe7] = 8'h00;
vram[12'hbe8] = 8'h70;
vram[12'hbe9] = 8'h18;
vram[12'hbea] = 8'h18;
vram[12'hbeb] = 8'h0e;
vram[12'hbec] = 8'h18;
vram[12'hbed] = 8'h18;
vram[12'hbee] = 8'h70;
vram[12'hbef] = 8'h00;
vram[12'hbf0] = 8'h76;
vram[12'hbf1] = 8'hdc;
vram[12'hbf2] = 8'h00;
vram[12'hbf3] = 8'h00;
vram[12'hbf4] = 8'h00;
vram[12'hbf5] = 8'h00;
vram[12'hbf6] = 8'h00;
vram[12'hbf7] = 8'h00;
vram[12'hbf8] = 8'hc0;
vram[12'hbf9] = 8'ha0;
vram[12'hbfa] = 8'hae;
vram[12'hbfb] = 8'ha4;
vram[12'hbfc] = 8'hc4;
vram[12'hbfd] = 8'h04;
vram[12'hbfe] = 8'h04;
vram[12'hbff] = 8'h00;
vram[12'hc00] = 8'h03;
vram[12'hc01] = 8'h03;
vram[12'hc02] = 8'h03;
vram[12'hc03] = 8'h03;
vram[12'hc04] = 8'h03;
vram[12'hc05] = 8'h03;
vram[12'hc06] = 8'h03;
vram[12'hc07] = 8'h03;
vram[12'hc08] = 8'h07;
vram[12'hc09] = 8'h07;
vram[12'hc0a] = 8'h07;
vram[12'hc0b] = 8'h07;
vram[12'hc0c] = 8'h07;
vram[12'hc0d] = 8'h07;
vram[12'hc0e] = 8'h07;
vram[12'hc0f] = 8'h07;
vram[12'hc10] = 8'h1f;
vram[12'hc11] = 8'h1f;
vram[12'hc12] = 8'h1f;
vram[12'hc13] = 8'h1f;
vram[12'hc14] = 8'h1f;
vram[12'hc15] = 8'h1f;
vram[12'hc16] = 8'h1f;
vram[12'hc17] = 8'h1f;
vram[12'hc18] = 8'h3f;
vram[12'hc19] = 8'h3f;
vram[12'hc1a] = 8'h3f;
vram[12'hc1b] = 8'h3f;
vram[12'hc1c] = 8'h3f;
vram[12'hc1d] = 8'h3f;
vram[12'hc1e] = 8'h3f;
vram[12'hc1f] = 8'h3f;
vram[12'hc20] = 8'h7f;
vram[12'hc21] = 8'h7f;
vram[12'hc22] = 8'h7f;
vram[12'hc23] = 8'h7f;
vram[12'hc24] = 8'h7f;
vram[12'hc25] = 8'h7f;
vram[12'hc26] = 8'h7f;
vram[12'hc27] = 8'h7f;
vram[12'hc28] = 8'hff;
vram[12'hc29] = 8'hff;
vram[12'hc2a] = 8'h00;
vram[12'hc2b] = 8'h00;
vram[12'hc2c] = 8'h00;
vram[12'hc2d] = 8'h00;
vram[12'hc2e] = 8'h00;
vram[12'hc2f] = 8'h00;
vram[12'hc30] = 8'hff;
vram[12'hc31] = 8'hff;
vram[12'hc32] = 8'hff;
vram[12'hc33] = 8'h00;
vram[12'hc34] = 8'h00;
vram[12'hc35] = 8'h00;
vram[12'hc36] = 8'h00;
vram[12'hc37] = 8'h00;
vram[12'hc38] = 8'hff;
vram[12'hc39] = 8'hff;
vram[12'hc3a] = 8'hff;
vram[12'hc3b] = 8'hff;
vram[12'hc3c] = 8'hff;
vram[12'hc3d] = 8'h00;
vram[12'hc3e] = 8'h00;
vram[12'hc3f] = 8'h00;
vram[12'hc40] = 8'hff;
vram[12'hc41] = 8'hff;
vram[12'hc42] = 8'hff;
vram[12'hc43] = 8'hff;
vram[12'hc44] = 8'hff;
vram[12'hc45] = 8'hff;
vram[12'hc46] = 8'h00;
vram[12'hc47] = 8'h00;
vram[12'hc48] = 8'hff;
vram[12'hc49] = 8'hff;
vram[12'hc4a] = 8'hff;
vram[12'hc4b] = 8'hff;
vram[12'hc4c] = 8'hff;
vram[12'hc4d] = 8'hff;
vram[12'hc4e] = 8'hff;
vram[12'hc4f] = 8'h00;
vram[12'hc50] = 8'haa;
vram[12'hc51] = 8'h55;
vram[12'hc52] = 8'haa;
vram[12'hc53] = 8'h55;
vram[12'hc54] = 8'h00;
vram[12'hc55] = 8'h00;
vram[12'hc56] = 8'h00;
vram[12'hc57] = 8'h00;
vram[12'hc58] = 8'h00;
vram[12'hc59] = 8'h00;
vram[12'hc5a] = 8'h00;
vram[12'hc5b] = 8'h00;
vram[12'hc5c] = 8'haa;
vram[12'hc5d] = 8'h55;
vram[12'hc5e] = 8'haa;
vram[12'hc5f] = 8'h55;
vram[12'hc60] = 8'ha0;
vram[12'hc61] = 8'h50;
vram[12'hc62] = 8'ha0;
vram[12'hc63] = 8'h50;
vram[12'hc64] = 8'ha0;
vram[12'hc65] = 8'h50;
vram[12'hc66] = 8'ha0;
vram[12'hc67] = 8'h50;
vram[12'hc68] = 8'h0a;
vram[12'hc69] = 8'h05;
vram[12'hc6a] = 8'h0a;
vram[12'hc6b] = 8'h05;
vram[12'hc6c] = 8'h0a;
vram[12'hc6d] = 8'h05;
vram[12'hc6e] = 8'h0a;
vram[12'hc6f] = 8'h05;
vram[12'hc70] = 8'hcc;
vram[12'hc71] = 8'hcc;
vram[12'hc72] = 8'h33;
vram[12'hc73] = 8'h33;
vram[12'hc74] = 8'h00;
vram[12'hc75] = 8'h00;
vram[12'hc76] = 8'h00;
vram[12'hc77] = 8'h00;
vram[12'hc78] = 8'h00;
vram[12'hc79] = 8'h00;
vram[12'hc7a] = 8'h00;
vram[12'hc7b] = 8'h00;
vram[12'hc7c] = 8'hcc;
vram[12'hc7d] = 8'hcc;
vram[12'hc7e] = 8'h33;
vram[12'hc7f] = 8'h33;
vram[12'hc80] = 8'hc0;
vram[12'hc81] = 8'hc0;
vram[12'hc82] = 8'h30;
vram[12'hc83] = 8'h30;
vram[12'hc84] = 8'hc0;
vram[12'hc85] = 8'hc0;
vram[12'hc86] = 8'h30;
vram[12'hc87] = 8'h30;
vram[12'hc88] = 8'h0c;
vram[12'hc89] = 8'h0c;
vram[12'hc8a] = 8'h03;
vram[12'hc8b] = 8'h03;
vram[12'hc8c] = 8'h0c;
vram[12'hc8d] = 8'h0c;
vram[12'hc8e] = 8'h03;
vram[12'hc8f] = 8'h03;
vram[12'hc90] = 8'h00;
vram[12'hc91] = 8'h01;
vram[12'hc92] = 8'h02;
vram[12'hc93] = 8'h05;
vram[12'hc94] = 8'h0a;
vram[12'hc95] = 8'h15;
vram[12'hc96] = 8'h2a;
vram[12'hc97] = 8'h55;
vram[12'hc98] = 8'h00;
vram[12'hc99] = 8'h80;
vram[12'hc9a] = 8'h40;
vram[12'hc9b] = 8'ha0;
vram[12'hc9c] = 8'h50;
vram[12'hc9d] = 8'ha8;
vram[12'hc9e] = 8'h54;
vram[12'hc9f] = 8'haa;
vram[12'hca0] = 8'haa;
vram[12'hca1] = 8'h54;
vram[12'hca2] = 8'ha8;
vram[12'hca3] = 8'h50;
vram[12'hca4] = 8'ha0;
vram[12'hca5] = 8'h40;
vram[12'hca6] = 8'h80;
vram[12'hca7] = 8'h00;
vram[12'hca8] = 8'haa;
vram[12'hca9] = 8'h55;
vram[12'hcaa] = 8'h2a;
vram[12'hcab] = 8'h15;
vram[12'hcac] = 8'h0a;
vram[12'hcad] = 8'h05;
vram[12'hcae] = 8'h02;
vram[12'hcaf] = 8'h01;
vram[12'hcb0] = 8'h00;
vram[12'hcb1] = 8'h00;
vram[12'hcb2] = 8'h01;
vram[12'hcb3] = 8'h03;
vram[12'hcb4] = 8'h0f;
vram[12'hcb5] = 8'h1f;
vram[12'hcb6] = 8'h3f;
vram[12'hcb7] = 8'h7f;
vram[12'hcb8] = 8'h00;
vram[12'hcb9] = 8'h00;
vram[12'hcba] = 8'h80;
vram[12'hcbb] = 8'hc0;
vram[12'hcbc] = 8'hf0;
vram[12'hcbd] = 8'hf8;
vram[12'hcbe] = 8'hfc;
vram[12'hcbf] = 8'hfe;
vram[12'hcc0] = 8'hfe;
vram[12'hcc1] = 8'hfc;
vram[12'hcc2] = 8'hf8;
vram[12'hcc3] = 8'hf0;
vram[12'hcc4] = 8'hc0;
vram[12'hcc5] = 8'h80;
vram[12'hcc6] = 8'h00;
vram[12'hcc7] = 8'h00;
vram[12'hcc8] = 8'h7f;
vram[12'hcc9] = 8'h3f;
vram[12'hcca] = 8'h1f;
vram[12'hccb] = 8'h0f;
vram[12'hccc] = 8'h03;
vram[12'hccd] = 8'h01;
vram[12'hcce] = 8'h00;
vram[12'hccf] = 8'h00;
vram[12'hcd0] = 8'hff;
vram[12'hcd1] = 8'hff;
vram[12'hcd2] = 8'hfe;
vram[12'hcd3] = 8'hfc;
vram[12'hcd4] = 8'hf0;
vram[12'hcd5] = 8'he0;
vram[12'hcd6] = 8'hc0;
vram[12'hcd7] = 8'h80;
vram[12'hcd8] = 8'hff;
vram[12'hcd9] = 8'hff;
vram[12'hcda] = 8'h7f;
vram[12'hcdb] = 8'h3f;
vram[12'hcdc] = 8'h0f;
vram[12'hcdd] = 8'h07;
vram[12'hcde] = 8'h03;
vram[12'hcdf] = 8'h01;
vram[12'hce0] = 8'h01;
vram[12'hce1] = 8'h03;
vram[12'hce2] = 8'h07;
vram[12'hce3] = 8'h0f;
vram[12'hce4] = 8'h3f;
vram[12'hce5] = 8'h7f;
vram[12'hce6] = 8'hff;
vram[12'hce7] = 8'hff;
vram[12'hce8] = 8'h80;
vram[12'hce9] = 8'hc0;
vram[12'hcea] = 8'he0;
vram[12'hceb] = 8'hf0;
vram[12'hcec] = 8'hfc;
vram[12'hced] = 8'hfe;
vram[12'hcee] = 8'hff;
vram[12'hcef] = 8'hff;
vram[12'hcf0] = 8'h00;
vram[12'hcf1] = 8'h00;
vram[12'hcf2] = 8'h00;
vram[12'hcf3] = 8'h00;
vram[12'hcf4] = 8'h03;
vram[12'hcf5] = 8'h0f;
vram[12'hcf6] = 8'h3f;
vram[12'hcf7] = 8'hff;
vram[12'hcf8] = 8'h00;
vram[12'hcf9] = 8'h00;
vram[12'hcfa] = 8'h00;
vram[12'hcfb] = 8'h00;
vram[12'hcfc] = 8'hc0;
vram[12'hcfd] = 8'hf0;
vram[12'hcfe] = 8'hfc;
vram[12'hcff] = 8'hff;
vram[12'hd00] = 8'hff;
vram[12'hd01] = 8'hfc;
vram[12'hd02] = 8'hf0;
vram[12'hd03] = 8'hc0;
vram[12'hd04] = 8'h00;
vram[12'hd05] = 8'h00;
vram[12'hd06] = 8'h00;
vram[12'hd07] = 8'h00;
vram[12'hd08] = 8'hff;
vram[12'hd09] = 8'h3f;
vram[12'hd0a] = 8'h0f;
vram[12'hd0b] = 8'h03;
vram[12'hd0c] = 8'h00;
vram[12'hd0d] = 8'h00;
vram[12'hd0e] = 8'h00;
vram[12'hd0f] = 8'h00;
vram[12'hd10] = 8'hff;
vram[12'hd11] = 8'hff;
vram[12'hd12] = 8'hff;
vram[12'hd13] = 8'hff;
vram[12'hd14] = 8'hfc;
vram[12'hd15] = 8'hf0;
vram[12'hd16] = 8'hc0;
vram[12'hd17] = 8'h00;
vram[12'hd18] = 8'hff;
vram[12'hd19] = 8'hff;
vram[12'hd1a] = 8'hff;
vram[12'hd1b] = 8'hff;
vram[12'hd1c] = 8'h3f;
vram[12'hd1d] = 8'h0f;
vram[12'hd1e] = 8'h03;
vram[12'hd1f] = 8'h00;
vram[12'hd20] = 8'h00;
vram[12'hd21] = 8'h03;
vram[12'hd22] = 8'h0f;
vram[12'hd23] = 8'h3f;
vram[12'hd24] = 8'hff;
vram[12'hd25] = 8'hff;
vram[12'hd26] = 8'hff;
vram[12'hd27] = 8'hff;
vram[12'hd28] = 8'h00;
vram[12'hd29] = 8'hc0;
vram[12'hd2a] = 8'hf0;
vram[12'hd2b] = 8'hfc;
vram[12'hd2c] = 8'hff;
vram[12'hd2d] = 8'hff;
vram[12'hd2e] = 8'hff;
vram[12'hd2f] = 8'hff;
vram[12'hd30] = 8'h01;
vram[12'hd31] = 8'h01;
vram[12'hd32] = 8'h03;
vram[12'hd33] = 8'h03;
vram[12'hd34] = 8'h07;
vram[12'hd35] = 8'h07;
vram[12'hd36] = 8'h0f;
vram[12'hd37] = 8'h0f;
vram[12'hd38] = 8'h80;
vram[12'hd39] = 8'h80;
vram[12'hd3a] = 8'hc0;
vram[12'hd3b] = 8'hc0;
vram[12'hd3c] = 8'he0;
vram[12'hd3d] = 8'he0;
vram[12'hd3e] = 8'hf0;
vram[12'hd3f] = 8'hf0;
vram[12'hd40] = 8'hf0;
vram[12'hd41] = 8'hf0;
vram[12'hd42] = 8'he0;
vram[12'hd43] = 8'he0;
vram[12'hd44] = 8'hc0;
vram[12'hd45] = 8'hc0;
vram[12'hd46] = 8'h80;
vram[12'hd47] = 8'h80;
vram[12'hd48] = 8'h0f;
vram[12'hd49] = 8'h0f;
vram[12'hd4a] = 8'h07;
vram[12'hd4b] = 8'h07;
vram[12'hd4c] = 8'h03;
vram[12'hd4d] = 8'h03;
vram[12'hd4e] = 8'h01;
vram[12'hd4f] = 8'h01;
vram[12'hd50] = 8'hfe;
vram[12'hd51] = 8'hfe;
vram[12'hd52] = 8'hfc;
vram[12'hd53] = 8'hfc;
vram[12'hd54] = 8'hf8;
vram[12'hd55] = 8'hf8;
vram[12'hd56] = 8'hf0;
vram[12'hd57] = 8'hf0;
vram[12'hd58] = 8'h7f;
vram[12'hd59] = 8'h7f;
vram[12'hd5a] = 8'h3f;
vram[12'hd5b] = 8'h3f;
vram[12'hd5c] = 8'h1f;
vram[12'hd5d] = 8'h1f;
vram[12'hd5e] = 8'h0f;
vram[12'hd5f] = 8'h0f;
vram[12'hd60] = 8'h0f;
vram[12'hd61] = 8'h0f;
vram[12'hd62] = 8'h1f;
vram[12'hd63] = 8'h1f;
vram[12'hd64] = 8'h3f;
vram[12'hd65] = 8'h3f;
vram[12'hd66] = 8'h7f;
vram[12'hd67] = 8'h7f;
vram[12'hd68] = 8'hf0;
vram[12'hd69] = 8'hf0;
vram[12'hd6a] = 8'hf8;
vram[12'hd6b] = 8'hf8;
vram[12'hd6c] = 8'hfc;
vram[12'hd6d] = 8'hfc;
vram[12'hd6e] = 8'hfe;
vram[12'hd6f] = 8'hfe;
vram[12'hd70] = 8'h00;
vram[12'hd71] = 8'h00;
vram[12'hd72] = 8'h00;
vram[12'hd73] = 8'h00;
vram[12'hd74] = 8'h00;
vram[12'hd75] = 8'h03;
vram[12'hd76] = 8'h1f;
vram[12'hd77] = 8'hff;
vram[12'hd78] = 8'h00;
vram[12'hd79] = 8'h00;
vram[12'hd7a] = 8'h00;
vram[12'hd7b] = 8'h00;
vram[12'hd7c] = 8'h00;
vram[12'hd7d] = 8'hc0;
vram[12'hd7e] = 8'hf8;
vram[12'hd7f] = 8'hff;
vram[12'hd80] = 8'hff;
vram[12'hd81] = 8'hf8;
vram[12'hd82] = 8'hc0;
vram[12'hd83] = 8'h00;
vram[12'hd84] = 8'h00;
vram[12'hd85] = 8'h00;
vram[12'hd86] = 8'h00;
vram[12'hd87] = 8'h00;
vram[12'hd88] = 8'hff;
vram[12'hd89] = 8'h1f;
vram[12'hd8a] = 8'h03;
vram[12'hd8b] = 8'h00;
vram[12'hd8c] = 8'h00;
vram[12'hd8d] = 8'h00;
vram[12'hd8e] = 8'h00;
vram[12'hd8f] = 8'h00;
vram[12'hd90] = 8'hff;
vram[12'hd91] = 8'hff;
vram[12'hd92] = 8'hff;
vram[12'hd93] = 8'hff;
vram[12'hd94] = 8'hff;
vram[12'hd95] = 8'hfc;
vram[12'hd96] = 8'he0;
vram[12'hd97] = 8'h00;
vram[12'hd98] = 8'hff;
vram[12'hd99] = 8'hff;
vram[12'hd9a] = 8'hff;
vram[12'hd9b] = 8'hff;
vram[12'hd9c] = 8'hff;
vram[12'hd9d] = 8'h3f;
vram[12'hd9e] = 8'h07;
vram[12'hd9f] = 8'h00;
vram[12'hda0] = 8'h00;
vram[12'hda1] = 8'h07;
vram[12'hda2] = 8'h3f;
vram[12'hda3] = 8'hff;
vram[12'hda4] = 8'hff;
vram[12'hda5] = 8'hff;
vram[12'hda6] = 8'hff;
vram[12'hda7] = 8'hff;
vram[12'hda8] = 8'h00;
vram[12'hda9] = 8'he0;
vram[12'hdaa] = 8'hfc;
vram[12'hdab] = 8'hff;
vram[12'hdac] = 8'hff;
vram[12'hdad] = 8'hff;
vram[12'hdae] = 8'hff;
vram[12'hdaf] = 8'hff;
vram[12'hdb0] = 8'h00;
vram[12'hdb1] = 8'h00;
vram[12'hdb2] = 8'h01;
vram[12'hdb3] = 8'h03;
vram[12'hdb4] = 8'h03;
vram[12'hdb5] = 8'h07;
vram[12'hdb6] = 8'h0f;
vram[12'hdb7] = 8'h0f;
vram[12'hdb8] = 8'h00;
vram[12'hdb9] = 8'h00;
vram[12'hdba] = 8'h80;
vram[12'hdbb] = 8'hc0;
vram[12'hdbc] = 8'hc0;
vram[12'hdbd] = 8'he0;
vram[12'hdbe] = 8'hf0;
vram[12'hdbf] = 8'hf0;
vram[12'hdc0] = 8'hf0;
vram[12'hdc1] = 8'hf0;
vram[12'hdc2] = 8'he0;
vram[12'hdc3] = 8'hc0;
vram[12'hdc4] = 8'hc0;
vram[12'hdc5] = 8'h80;
vram[12'hdc6] = 8'h00;
vram[12'hdc7] = 8'h00;
vram[12'hdc8] = 8'h0f;
vram[12'hdc9] = 8'h0f;
vram[12'hdca] = 8'h07;
vram[12'hdcb] = 8'h03;
vram[12'hdcc] = 8'h03;
vram[12'hdcd] = 8'h01;
vram[12'hdce] = 8'h00;
vram[12'hdcf] = 8'h00;
vram[12'hdd0] = 8'hff;
vram[12'hdd1] = 8'hff;
vram[12'hdd2] = 8'hfe;
vram[12'hdd3] = 8'hfc;
vram[12'hdd4] = 8'hfc;
vram[12'hdd5] = 8'hf8;
vram[12'hdd6] = 8'hf0;
vram[12'hdd7] = 8'hf0;
vram[12'hdd8] = 8'hff;
vram[12'hdd9] = 8'hff;
vram[12'hdda] = 8'h7f;
vram[12'hddb] = 8'h3f;
vram[12'hddc] = 8'h3f;
vram[12'hddd] = 8'h1f;
vram[12'hdde] = 8'h0f;
vram[12'hddf] = 8'h0f;
vram[12'hde0] = 8'h0f;
vram[12'hde1] = 8'h0f;
vram[12'hde2] = 8'h1f;
vram[12'hde3] = 8'h3f;
vram[12'hde4] = 8'h3f;
vram[12'hde5] = 8'h7f;
vram[12'hde6] = 8'hff;
vram[12'hde7] = 8'hff;
vram[12'hde8] = 8'hf0;
vram[12'hde9] = 8'hf0;
vram[12'hdea] = 8'hf8;
vram[12'hdeb] = 8'hfc;
vram[12'hdec] = 8'hfc;
vram[12'hded] = 8'hfe;
vram[12'hdee] = 8'hff;
vram[12'hdef] = 8'hff;
vram[12'hdf0] = 8'h00;
vram[12'hdf1] = 8'h00;
vram[12'hdf2] = 8'h00;
vram[12'hdf3] = 8'h00;
vram[12'hdf4] = 8'h01;
vram[12'hdf5] = 8'h03;
vram[12'hdf6] = 8'h07;
vram[12'hdf7] = 8'h0f;
vram[12'hdf8] = 8'h00;
vram[12'hdf9] = 8'h00;
vram[12'hdfa] = 8'h00;
vram[12'hdfb] = 8'h00;
vram[12'hdfc] = 8'h80;
vram[12'hdfd] = 8'hc0;
vram[12'hdfe] = 8'he0;
vram[12'hdff] = 8'hf0;
vram[12'he00] = 8'hf0;
vram[12'he01] = 8'he0;
vram[12'he02] = 8'hc0;
vram[12'he03] = 8'h80;
vram[12'he04] = 8'h00;
vram[12'he05] = 8'h00;
vram[12'he06] = 8'h00;
vram[12'he07] = 8'h00;
vram[12'he08] = 8'h0f;
vram[12'he09] = 8'h07;
vram[12'he0a] = 8'h03;
vram[12'he0b] = 8'h01;
vram[12'he0c] = 8'h00;
vram[12'he0d] = 8'h00;
vram[12'he0e] = 8'h00;
vram[12'he0f] = 8'h00;
vram[12'he10] = 8'hff;
vram[12'he11] = 8'hff;
vram[12'he12] = 8'hff;
vram[12'he13] = 8'hff;
vram[12'he14] = 8'hfe;
vram[12'he15] = 8'hfc;
vram[12'he16] = 8'hf8;
vram[12'he17] = 8'hf0;
vram[12'he18] = 8'hff;
vram[12'he19] = 8'hff;
vram[12'he1a] = 8'hff;
vram[12'he1b] = 8'hff;
vram[12'he1c] = 8'h7f;
vram[12'he1d] = 8'h3f;
vram[12'he1e] = 8'h1f;
vram[12'he1f] = 8'h0f;
vram[12'he20] = 8'h0f;
vram[12'he21] = 8'h1f;
vram[12'he22] = 8'h3f;
vram[12'he23] = 8'h7f;
vram[12'he24] = 8'hff;
vram[12'he25] = 8'hff;
vram[12'he26] = 8'hff;
vram[12'he27] = 8'hff;
vram[12'he28] = 8'hf0;
vram[12'he29] = 8'hf8;
vram[12'he2a] = 8'hfc;
vram[12'he2b] = 8'hfe;
vram[12'he2c] = 8'hff;
vram[12'he2d] = 8'hff;
vram[12'he2e] = 8'hff;
vram[12'he2f] = 8'hff;
vram[12'he30] = 8'h00;
vram[12'he31] = 8'h00;
vram[12'he32] = 8'h00;
vram[12'he33] = 8'h00;
vram[12'he34] = 8'h03;
vram[12'he35] = 8'h07;
vram[12'he36] = 8'h0f;
vram[12'he37] = 8'h0f;
vram[12'he38] = 8'h00;
vram[12'he39] = 8'h00;
vram[12'he3a] = 8'h00;
vram[12'he3b] = 8'h00;
vram[12'he3c] = 8'hc0;
vram[12'he3d] = 8'he0;
vram[12'he3e] = 8'hf0;
vram[12'he3f] = 8'hf0;
vram[12'he40] = 8'hf0;
vram[12'he41] = 8'hf0;
vram[12'he42] = 8'he0;
vram[12'he43] = 8'hc0;
vram[12'he44] = 8'h00;
vram[12'he45] = 8'h00;
vram[12'he46] = 8'h00;
vram[12'he47] = 8'h00;
vram[12'he48] = 8'h0f;
vram[12'he49] = 8'h0f;
vram[12'he4a] = 8'h07;
vram[12'he4b] = 8'h03;
vram[12'he4c] = 8'h00;
vram[12'he4d] = 8'h00;
vram[12'he4e] = 8'h00;
vram[12'he4f] = 8'h00;
vram[12'he50] = 8'h00;
vram[12'he51] = 8'h00;
vram[12'he52] = 8'h00;
vram[12'he53] = 8'h00;
vram[12'he54] = 8'h00;
vram[12'he55] = 8'h01;
vram[12'he56] = 8'h03;
vram[12'he57] = 8'h07;
vram[12'he58] = 8'h00;
vram[12'he59] = 8'h00;
vram[12'he5a] = 8'h00;
vram[12'he5b] = 8'h00;
vram[12'he5c] = 8'h00;
vram[12'he5d] = 8'h80;
vram[12'he5e] = 8'hc0;
vram[12'he5f] = 8'he0;
vram[12'he60] = 8'he0;
vram[12'he61] = 8'hc0;
vram[12'he62] = 8'h80;
vram[12'he63] = 8'h00;
vram[12'he64] = 8'h00;
vram[12'he65] = 8'h00;
vram[12'he66] = 8'h00;
vram[12'he67] = 8'h00;
vram[12'he68] = 8'h07;
vram[12'he69] = 8'h03;
vram[12'he6a] = 8'h01;
vram[12'he6b] = 8'h00;
vram[12'he6c] = 8'h00;
vram[12'he6d] = 8'h00;
vram[12'he6e] = 8'h00;
vram[12'he6f] = 8'h00;
vram[12'he70] = 8'hff;
vram[12'he71] = 8'hff;
vram[12'he72] = 8'hff;
vram[12'he73] = 8'hff;
vram[12'he74] = 8'hff;
vram[12'he75] = 8'hfe;
vram[12'he76] = 8'hfc;
vram[12'he77] = 8'hf8;
vram[12'he78] = 8'hff;
vram[12'he79] = 8'hff;
vram[12'he7a] = 8'hff;
vram[12'he7b] = 8'hff;
vram[12'he7c] = 8'hff;
vram[12'he7d] = 8'h7f;
vram[12'he7e] = 8'h3f;
vram[12'he7f] = 8'h1f;
vram[12'he80] = 8'h1f;
vram[12'he81] = 8'h3f;
vram[12'he82] = 8'h7f;
vram[12'he83] = 8'hff;
vram[12'he84] = 8'hff;
vram[12'he85] = 8'hff;
vram[12'he86] = 8'hff;
vram[12'he87] = 8'hff;
vram[12'he88] = 8'hf8;
vram[12'he89] = 8'hfc;
vram[12'he8a] = 8'hfe;
vram[12'he8b] = 8'hff;
vram[12'he8c] = 8'hff;
vram[12'he8d] = 8'hff;
vram[12'he8e] = 8'hff;
vram[12'he8f] = 8'hff;
vram[12'he90] = 8'h00;
vram[12'he91] = 8'h00;
vram[12'he92] = 8'h00;
vram[12'he93] = 8'h03;
vram[12'he94] = 8'h3f;
vram[12'he95] = 8'hff;
vram[12'he96] = 8'hff;
vram[12'he97] = 8'hff;
vram[12'he98] = 8'h00;
vram[12'he99] = 8'h00;
vram[12'he9a] = 8'h00;
vram[12'he9b] = 8'hc0;
vram[12'he9c] = 8'hfc;
vram[12'he9d] = 8'hff;
vram[12'he9e] = 8'hff;
vram[12'he9f] = 8'hff;
vram[12'hea0] = 8'hff;
vram[12'hea1] = 8'hff;
vram[12'hea2] = 8'hff;
vram[12'hea3] = 8'hfc;
vram[12'hea4] = 8'hc0;
vram[12'hea5] = 8'h00;
vram[12'hea6] = 8'h00;
vram[12'hea7] = 8'h00;
vram[12'hea8] = 8'hff;
vram[12'hea9] = 8'hff;
vram[12'heaa] = 8'hff;
vram[12'heab] = 8'h3f;
vram[12'heac] = 8'h03;
vram[12'head] = 8'h00;
vram[12'heae] = 8'h00;
vram[12'heaf] = 8'h00;
vram[12'heb0] = 8'hef;
vram[12'heb1] = 8'hef;
vram[12'heb2] = 8'hc7;
vram[12'heb3] = 8'hc7;
vram[12'heb4] = 8'h83;
vram[12'heb5] = 8'h83;
vram[12'heb6] = 8'h01;
vram[12'heb7] = 8'h01;
vram[12'heb8] = 8'h3f;
vram[12'heb9] = 8'h0f;
vram[12'heba] = 8'h03;
vram[12'hebb] = 8'h00;
vram[12'hebc] = 8'h03;
vram[12'hebd] = 8'h0f;
vram[12'hebe] = 8'h3f;
vram[12'hebf] = 8'hff;
vram[12'hec0] = 8'h01;
vram[12'hec1] = 8'h01;
vram[12'hec2] = 8'h83;
vram[12'hec3] = 8'h83;
vram[12'hec4] = 8'hc7;
vram[12'hec5] = 8'hc7;
vram[12'hec6] = 8'hef;
vram[12'hec7] = 8'hef;
vram[12'hec8] = 8'hfc;
vram[12'hec9] = 8'hf0;
vram[12'heca] = 8'hc0;
vram[12'hecb] = 8'h00;
vram[12'hecc] = 8'hc0;
vram[12'hecd] = 8'hf0;
vram[12'hece] = 8'hfc;
vram[12'hecf] = 8'hff;
vram[12'hed0] = 8'h00;
vram[12'hed1] = 8'h00;
vram[12'hed2] = 8'h00;
vram[12'hed3] = 8'h00;
vram[12'hed4] = 8'h10;
vram[12'hed5] = 8'h38;
vram[12'hed6] = 8'h7c;
vram[12'hed7] = 8'hfe;
vram[12'hed8] = 8'h80;
vram[12'hed9] = 8'hc0;
vram[12'heda] = 8'he0;
vram[12'hedb] = 8'hf0;
vram[12'hedc] = 8'he0;
vram[12'hedd] = 8'hc0;
vram[12'hede] = 8'h80;
vram[12'hedf] = 8'h00;
vram[12'hee0] = 8'hfe;
vram[12'hee1] = 8'h7c;
vram[12'hee2] = 8'h38;
vram[12'hee3] = 8'h10;
vram[12'hee4] = 8'h00;
vram[12'hee5] = 8'h00;
vram[12'hee6] = 8'h00;
vram[12'hee7] = 8'h00;
vram[12'hee8] = 8'h01;
vram[12'hee9] = 8'h03;
vram[12'heea] = 8'h07;
vram[12'heeb] = 8'h0f;
vram[12'heec] = 8'h07;
vram[12'heed] = 8'h03;
vram[12'heee] = 8'h01;
vram[12'heef] = 8'h00;
vram[12'hef0] = 8'hff;
vram[12'hef1] = 8'hff;
vram[12'hef2] = 8'hff;
vram[12'hef3] = 8'hff;
vram[12'hef4] = 8'hef;
vram[12'hef5] = 8'hc7;
vram[12'hef6] = 8'h83;
vram[12'hef7] = 8'h01;
vram[12'hef8] = 8'h7f;
vram[12'hef9] = 8'h3f;
vram[12'hefa] = 8'h1f;
vram[12'hefb] = 8'h0f;
vram[12'hefc] = 8'h1f;
vram[12'hefd] = 8'h3f;
vram[12'hefe] = 8'h7f;
vram[12'heff] = 8'hff;
vram[12'hf00] = 8'h01;
vram[12'hf01] = 8'h83;
vram[12'hf02] = 8'hc7;
vram[12'hf03] = 8'hef;
vram[12'hf04] = 8'hff;
vram[12'hf05] = 8'hff;
vram[12'hf06] = 8'hff;
vram[12'hf07] = 8'hff;
vram[12'hf08] = 8'hfe;
vram[12'hf09] = 8'hfc;
vram[12'hf0a] = 8'hf8;
vram[12'hf0b] = 8'hf0;
vram[12'hf0c] = 8'hf8;
vram[12'hf0d] = 8'hfc;
vram[12'hf0e] = 8'hfe;
vram[12'hf0f] = 8'hff;
vram[12'hf10] = 8'h18;
vram[12'hf11] = 8'h3c;
vram[12'hf12] = 8'h7e;
vram[12'hf13] = 8'hff;
vram[12'hf14] = 8'hff;
vram[12'hf15] = 8'hff;
vram[12'hf16] = 8'hff;
vram[12'hf17] = 8'hff;
vram[12'hf18] = 8'hf8;
vram[12'hf19] = 8'hfc;
vram[12'hf1a] = 8'hfe;
vram[12'hf1b] = 8'hff;
vram[12'hf1c] = 8'hff;
vram[12'hf1d] = 8'hfe;
vram[12'hf1e] = 8'hfc;
vram[12'hf1f] = 8'hf8;
vram[12'hf20] = 8'hff;
vram[12'hf21] = 8'hff;
vram[12'hf22] = 8'hff;
vram[12'hf23] = 8'hff;
vram[12'hf24] = 8'hff;
vram[12'hf25] = 8'h7e;
vram[12'hf26] = 8'h3c;
vram[12'hf27] = 8'h18;
vram[12'hf28] = 8'h1f;
vram[12'hf29] = 8'h3f;
vram[12'hf2a] = 8'h7f;
vram[12'hf2b] = 8'hff;
vram[12'hf2c] = 8'hff;
vram[12'hf2d] = 8'h7f;
vram[12'hf2e] = 8'h3f;
vram[12'hf2f] = 8'h1f;
vram[12'hf30] = 8'he7;
vram[12'hf31] = 8'hc3;
vram[12'hf32] = 8'h81;
vram[12'hf33] = 8'h00;
vram[12'hf34] = 8'h00;
vram[12'hf35] = 8'h00;
vram[12'hf36] = 8'h00;
vram[12'hf37] = 8'h00;
vram[12'hf38] = 8'h07;
vram[12'hf39] = 8'h03;
vram[12'hf3a] = 8'h01;
vram[12'hf3b] = 8'h00;
vram[12'hf3c] = 8'h00;
vram[12'hf3d] = 8'h01;
vram[12'hf3e] = 8'h03;
vram[12'hf3f] = 8'h07;
vram[12'hf40] = 8'h00;
vram[12'hf41] = 8'h00;
vram[12'hf42] = 8'h00;
vram[12'hf43] = 8'h00;
vram[12'hf44] = 8'h00;
vram[12'hf45] = 8'h81;
vram[12'hf46] = 8'hc3;
vram[12'hf47] = 8'he7;
vram[12'hf48] = 8'he0;
vram[12'hf49] = 8'hc0;
vram[12'hf4a] = 8'h80;
vram[12'hf4b] = 8'h00;
vram[12'hf4c] = 8'h00;
vram[12'hf4d] = 8'h80;
vram[12'hf4e] = 8'hc0;
vram[12'hf4f] = 8'he0;
vram[12'hf50] = 8'hff;
vram[12'hf51] = 8'h7e;
vram[12'hf52] = 8'h3c;
vram[12'hf53] = 8'h18;
vram[12'hf54] = 8'h18;
vram[12'hf55] = 8'h3c;
vram[12'hf56] = 8'h7e;
vram[12'hf57] = 8'hff;
vram[12'hf58] = 8'h81;
vram[12'hf59] = 8'hc3;
vram[12'hf5a] = 8'he7;
vram[12'hf5b] = 8'hff;
vram[12'hf5c] = 8'hff;
vram[12'hf5d] = 8'he7;
vram[12'hf5e] = 8'hc3;
vram[12'hf5f] = 8'h81;
vram[12'hf60] = 8'hff;
vram[12'hf61] = 8'hff;
vram[12'hf62] = 8'hc0;
vram[12'hf63] = 8'hc0;
vram[12'hf64] = 8'hc0;
vram[12'hf65] = 8'hc0;
vram[12'hf66] = 8'hc0;
vram[12'hf67] = 8'hc0;
vram[12'hf68] = 8'hff;
vram[12'hf69] = 8'hff;
vram[12'hf6a] = 8'h03;
vram[12'hf6b] = 8'h03;
vram[12'hf6c] = 8'h03;
vram[12'hf6d] = 8'h03;
vram[12'hf6e] = 8'h03;
vram[12'hf6f] = 8'h03;
vram[12'hf70] = 8'h03;
vram[12'hf71] = 8'h03;
vram[12'hf72] = 8'h03;
vram[12'hf73] = 8'h03;
vram[12'hf74] = 8'h03;
vram[12'hf75] = 8'h03;
vram[12'hf76] = 8'hff;
vram[12'hf77] = 8'hff;
vram[12'hf78] = 8'hc0;
vram[12'hf79] = 8'hc0;
vram[12'hf7a] = 8'hc0;
vram[12'hf7b] = 8'hc0;
vram[12'hf7c] = 8'hc0;
vram[12'hf7d] = 8'hc0;
vram[12'hf7e] = 8'hff;
vram[12'hf7f] = 8'hff;
vram[12'hf80] = 8'h00;
vram[12'hf81] = 8'hff;
vram[12'hf82] = 8'hff;
vram[12'hf83] = 8'h00;
vram[12'hf84] = 8'h00;
vram[12'hf85] = 8'h00;
vram[12'hf86] = 8'h00;
vram[12'hf87] = 8'h00;
vram[12'hf88] = 8'h00;
vram[12'hf89] = 8'h00;
vram[12'hf8a] = 8'hff;
vram[12'hf8b] = 8'hff;
vram[12'hf8c] = 8'h00;
vram[12'hf8d] = 8'h00;
vram[12'hf8e] = 8'h00;
vram[12'hf8f] = 8'h00;
vram[12'hf90] = 8'h00;
vram[12'hf91] = 8'h00;
vram[12'hf92] = 8'h00;
vram[12'hf93] = 8'hff;
vram[12'hf94] = 8'hff;
vram[12'hf95] = 8'h00;
vram[12'hf96] = 8'h00;
vram[12'hf97] = 8'h00;
vram[12'hf98] = 8'h00;
vram[12'hf99] = 8'h00;
vram[12'hf9a] = 8'h00;
vram[12'hf9b] = 8'h00;
vram[12'hf9c] = 8'hff;
vram[12'hf9d] = 8'hff;
vram[12'hf9e] = 8'h00;
vram[12'hf9f] = 8'h00;
vram[12'hfa0] = 8'h00;
vram[12'hfa1] = 8'h00;
vram[12'hfa2] = 8'h00;
vram[12'hfa3] = 8'h00;
vram[12'hfa4] = 8'h00;
vram[12'hfa5] = 8'hff;
vram[12'hfa6] = 8'hff;
vram[12'hfa7] = 8'h00;
vram[12'hfa8] = 8'h60;
vram[12'hfa9] = 8'h60;
vram[12'hfaa] = 8'h60;
vram[12'hfab] = 8'h60;
vram[12'hfac] = 8'h60;
vram[12'hfad] = 8'h60;
vram[12'hfae] = 8'h60;
vram[12'hfaf] = 8'h60;
vram[12'hfb0] = 8'h30;
vram[12'hfb1] = 8'h30;
vram[12'hfb2] = 8'h30;
vram[12'hfb3] = 8'h30;
vram[12'hfb4] = 8'h30;
vram[12'hfb5] = 8'h30;
vram[12'hfb6] = 8'h30;
vram[12'hfb7] = 8'h30;
vram[12'hfb8] = 8'h0c;
vram[12'hfb9] = 8'h0c;
vram[12'hfba] = 8'h0c;
vram[12'hfbb] = 8'h0c;
vram[12'hfbc] = 8'h0c;
vram[12'hfbd] = 8'h0c;
vram[12'hfbe] = 8'h0c;
vram[12'hfbf] = 8'h0c;
vram[12'hfc0] = 8'h06;
vram[12'hfc1] = 8'h06;
vram[12'hfc2] = 8'h06;
vram[12'hfc3] = 8'h06;
vram[12'hfc4] = 8'h06;
vram[12'hfc5] = 8'h06;
vram[12'hfc6] = 8'h06;
vram[12'hfc7] = 8'h06;
vram[12'hfc8] = 8'he0;
vram[12'hfc9] = 8'h38;
vram[12'hfca] = 8'h0e;
vram[12'hfcb] = 8'h03;
vram[12'hfcc] = 8'h00;
vram[12'hfcd] = 8'h00;
vram[12'hfce] = 8'h00;
vram[12'hfcf] = 8'h00;
vram[12'hfd0] = 8'h00;
vram[12'hfd1] = 8'h00;
vram[12'hfd2] = 8'h00;
vram[12'hfd3] = 8'h80;
vram[12'hfd4] = 8'he0;
vram[12'hfd5] = 8'h38;
vram[12'hfd6] = 8'h0e;
vram[12'hfd7] = 8'h03;
vram[12'hfd8] = 8'h00;
vram[12'hfd9] = 8'h00;
vram[12'hfda] = 8'h00;
vram[12'hfdb] = 8'h01;
vram[12'hfdc] = 8'h07;
vram[12'hfdd] = 8'h1c;
vram[12'hfde] = 8'h70;
vram[12'hfdf] = 8'hc0;
vram[12'hfe0] = 8'h07;
vram[12'hfe1] = 8'h1c;
vram[12'hfe2] = 8'h70;
vram[12'hfe3] = 8'hc0;
vram[12'hfe4] = 8'h00;
vram[12'hfe5] = 8'h00;
vram[12'hfe6] = 8'h00;
vram[12'hfe7] = 8'h00;
vram[12'hfe8] = 8'h80;
vram[12'hfe9] = 8'hc0;
vram[12'hfea] = 8'hc0;
vram[12'hfeb] = 8'h60;
vram[12'hfec] = 8'h60;
vram[12'hfed] = 8'h30;
vram[12'hfee] = 8'h30;
vram[12'hfef] = 8'h18;
vram[12'hff0] = 8'h18;
vram[12'hff1] = 8'h0c;
vram[12'hff2] = 8'h0c;
vram[12'hff3] = 8'h06;
vram[12'hff4] = 8'h06;
vram[12'hff5] = 8'h03;
vram[12'hff6] = 8'h03;
vram[12'hff7] = 8'h01;
vram[12'hff8] = 8'h18;
vram[12'hff9] = 8'h30;
vram[12'hffa] = 8'h30;
vram[12'hffb] = 8'h60;
vram[12'hffc] = 8'h60;
vram[12'hffd] = 8'hc0;
vram[12'hffe] = 8'hc0;
vram[12'hfff] = 8'h80;
