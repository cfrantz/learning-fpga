mem[0] = 8'h1c;
mem[1] = 8'h1d;
mem[2] = 8'h1c;
mem[3] = 8'h1d;
mem[4] = 8'h1c;
mem[5] = 8'h1d;
mem[6] = 8'h1c;
mem[7] = 8'h1d;
mem[8] = 8'h1c;
mem[9] = 8'h1d;
mem[10] = 8'h1c;
mem[11] = 8'h1d;
mem[12] = 8'h1c;
mem[13] = 8'h1d;
mem[14] = 8'h1c;
mem[15] = 8'h1d;
mem[16] = 8'h1c;
mem[17] = 8'h1d;
mem[18] = 8'h1c;
mem[19] = 8'h1d;
mem[20] = 8'h1c;
mem[21] = 8'h1d;
mem[22] = 8'h1c;
mem[23] = 8'h1d;
mem[24] = 8'h1c;
mem[25] = 8'h1d;
mem[26] = 8'h1c;
mem[27] = 8'h1d;
mem[28] = 8'h1c;
mem[29] = 8'h1d;
mem[30] = 8'h1c;
mem[31] = 8'h1d;
mem[32] = 8'h20;
mem[33] = 8'h20;
mem[34] = 8'h20;
mem[35] = 8'h20;
mem[36] = 8'h20;
mem[37] = 8'h20;
mem[38] = 8'h20;
mem[39] = 8'h20;
mem[40] = 8'h20;
mem[41] = 8'h20;
mem[42] = 8'h20;
mem[43] = 8'h20;
mem[44] = 8'h20;
mem[45] = 8'h20;
mem[46] = 8'h20;
mem[47] = 8'h20;
mem[48] = 8'h20;
mem[49] = 8'h20;
mem[50] = 8'h20;
mem[51] = 8'h20;
mem[52] = 8'h20;
mem[53] = 8'h20;
mem[54] = 8'h20;
mem[55] = 8'h20;
mem[56] = 8'h20;
mem[57] = 8'h20;
mem[58] = 8'h20;
mem[59] = 8'h20;
mem[60] = 8'h20;
mem[61] = 8'h20;
mem[62] = 8'h20;
mem[63] = 8'h20;
mem[64] = 8'h54;
mem[65] = 8'h69;
mem[66] = 8'h6e;
mem[67] = 8'h79;
mem[68] = 8'h36;
mem[69] = 8'h35;
mem[70] = 8'h30;
mem[71] = 8'h32;
mem[72] = 8'h20;
mem[73] = 8'h61;
mem[74] = 8'h6e;
mem[75] = 8'h64;
mem[76] = 8'h20;
mem[77] = 8'h54;
mem[78] = 8'h69;
mem[79] = 8'h6e;
mem[80] = 8'h79;
mem[81] = 8'h56;
mem[82] = 8'h47;
mem[83] = 8'h41;
mem[84] = 8'h20;
mem[85] = 8'h44;
mem[86] = 8'h69;
mem[87] = 8'h73;
mem[88] = 8'h70;
mem[89] = 8'h6c;
mem[90] = 8'h61;
mem[91] = 8'h79;
mem[92] = 8'h20;
mem[93] = 8'h20;
mem[94] = 8'h20;
mem[95] = 8'h20;
mem[96] = 8'h62;
mem[97] = 8'h79;
mem[98] = 8'h20;
mem[99] = 8'h43;
mem[100] = 8'h46;
mem[101] = 8'h32;
mem[102] = 8'h30;
mem[103] = 8'h37;
mem[104] = 8'h2e;
mem[105] = 8'h20;
mem[106] = 8'h20;
mem[107] = 8'h20;
mem[108] = 8'h20;
mem[109] = 8'h20;
mem[110] = 8'h20;
mem[111] = 8'h20;
mem[112] = 8'h20;
mem[113] = 8'h20;
mem[114] = 8'h20;
mem[115] = 8'h20;
mem[116] = 8'h20;
mem[117] = 8'h20;
mem[118] = 8'h20;
mem[119] = 8'h20;
mem[120] = 8'h20;
mem[121] = 8'h20;
mem[122] = 8'h20;
mem[123] = 8'h20;
mem[124] = 8'h20;
mem[125] = 8'h20;
mem[126] = 8'h20;
mem[127] = 8'h20;
mem[128] = 8'h00;
mem[129] = 8'h00;
mem[130] = 8'h00;
mem[131] = 8'h00;
mem[132] = 8'h00;
mem[133] = 8'h00;
mem[134] = 8'h00;
mem[135] = 8'h00;
mem[136] = 8'h00;
mem[137] = 8'h00;
mem[138] = 8'h00;
mem[139] = 8'h00;
mem[140] = 8'h00;
mem[141] = 8'h00;
mem[142] = 8'h00;
mem[143] = 8'h00;
mem[144] = 8'h00;
mem[145] = 8'h00;
mem[146] = 8'h00;
mem[147] = 8'h00;
mem[148] = 8'h00;
mem[149] = 8'h00;
mem[150] = 8'h00;
mem[151] = 8'h00;
mem[152] = 8'h00;
mem[153] = 8'h00;
mem[154] = 8'h00;
mem[155] = 8'h00;
mem[156] = 8'h00;
mem[157] = 8'h00;
mem[158] = 8'h00;
mem[159] = 8'h00;
mem[160] = 8'h00;
mem[161] = 8'h00;
mem[162] = 8'h00;
mem[163] = 8'h00;
mem[164] = 8'h00;
mem[165] = 8'h00;
mem[166] = 8'h00;
mem[167] = 8'h00;
mem[168] = 8'h00;
mem[169] = 8'h00;
mem[170] = 8'h00;
mem[171] = 8'h00;
mem[172] = 8'h00;
mem[173] = 8'h00;
mem[174] = 8'h00;
mem[175] = 8'h00;
mem[176] = 8'h00;
mem[177] = 8'h00;
mem[178] = 8'h00;
mem[179] = 8'h00;
mem[180] = 8'h00;
mem[181] = 8'h00;
mem[182] = 8'h00;
mem[183] = 8'h00;
mem[184] = 8'h00;
mem[185] = 8'h00;
mem[186] = 8'h00;
mem[187] = 8'h00;
mem[188] = 8'h00;
mem[189] = 8'h00;
mem[190] = 8'h00;
mem[191] = 8'h00;
mem[192] = 8'h00;
mem[193] = 8'h00;
mem[194] = 8'h00;
mem[195] = 8'h00;
mem[196] = 8'h00;
mem[197] = 8'h00;
mem[198] = 8'h00;
mem[199] = 8'h00;
mem[200] = 8'h00;
mem[201] = 8'h00;
mem[202] = 8'h00;
mem[203] = 8'h00;
mem[204] = 8'h00;
mem[205] = 8'h00;
mem[206] = 8'h00;
mem[207] = 8'h00;
mem[208] = 8'h00;
mem[209] = 8'h00;
mem[210] = 8'h00;
mem[211] = 8'h00;
mem[212] = 8'h00;
mem[213] = 8'h00;
mem[214] = 8'h00;
mem[215] = 8'h00;
mem[216] = 8'h00;
mem[217] = 8'h00;
mem[218] = 8'h00;
mem[219] = 8'h00;
mem[220] = 8'h00;
mem[221] = 8'h00;
mem[222] = 8'h00;
mem[223] = 8'h00;
mem[224] = 8'h00;
mem[225] = 8'h00;
mem[226] = 8'h00;
mem[227] = 8'h00;
mem[228] = 8'h00;
mem[229] = 8'h00;
mem[230] = 8'h00;
mem[231] = 8'h00;
mem[232] = 8'h00;
mem[233] = 8'h00;
mem[234] = 8'h00;
mem[235] = 8'h00;
mem[236] = 8'h00;
mem[237] = 8'h00;
mem[238] = 8'h00;
mem[239] = 8'h00;
mem[240] = 8'h00;
mem[241] = 8'h00;
mem[242] = 8'h00;
mem[243] = 8'h00;
mem[244] = 8'h00;
mem[245] = 8'h00;
mem[246] = 8'h00;
mem[247] = 8'h00;
mem[248] = 8'h00;
mem[249] = 8'h00;
mem[250] = 8'h00;
mem[251] = 8'h00;
mem[252] = 8'h00;
mem[253] = 8'h00;
mem[254] = 8'h00;
mem[255] = 8'h00;
mem[256] = 8'h00;
mem[257] = 8'h00;
mem[258] = 8'h00;
mem[259] = 8'h00;
mem[260] = 8'h00;
mem[261] = 8'h00;
mem[262] = 8'h00;
mem[263] = 8'h00;
mem[264] = 8'h00;
mem[265] = 8'h00;
mem[266] = 8'h00;
mem[267] = 8'h00;
mem[268] = 8'h00;
mem[269] = 8'h00;
mem[270] = 8'h00;
mem[271] = 8'h00;
mem[272] = 8'h00;
mem[273] = 8'h00;
mem[274] = 8'h00;
mem[275] = 8'h00;
mem[276] = 8'h00;
mem[277] = 8'h00;
mem[278] = 8'h00;
mem[279] = 8'h00;
mem[280] = 8'h00;
mem[281] = 8'h00;
mem[282] = 8'h00;
mem[283] = 8'h00;
mem[284] = 8'h00;
mem[285] = 8'h00;
mem[286] = 8'h00;
mem[287] = 8'h00;
mem[288] = 8'h00;
mem[289] = 8'h00;
mem[290] = 8'h00;
mem[291] = 8'h00;
mem[292] = 8'h00;
mem[293] = 8'h00;
mem[294] = 8'h00;
mem[295] = 8'h00;
mem[296] = 8'h00;
mem[297] = 8'h00;
mem[298] = 8'h00;
mem[299] = 8'h00;
mem[300] = 8'h00;
mem[301] = 8'h00;
mem[302] = 8'h00;
mem[303] = 8'h00;
mem[304] = 8'h00;
mem[305] = 8'h00;
mem[306] = 8'h00;
mem[307] = 8'h00;
mem[308] = 8'h00;
mem[309] = 8'h00;
mem[310] = 8'h00;
mem[311] = 8'h00;
mem[312] = 8'h00;
mem[313] = 8'h00;
mem[314] = 8'h00;
mem[315] = 8'h00;
mem[316] = 8'h00;
mem[317] = 8'h00;
mem[318] = 8'h00;
mem[319] = 8'h00;
mem[320] = 8'h00;
mem[321] = 8'h00;
mem[322] = 8'h00;
mem[323] = 8'h00;
mem[324] = 8'h00;
mem[325] = 8'h00;
mem[326] = 8'h00;
mem[327] = 8'h00;
mem[328] = 8'h00;
mem[329] = 8'h00;
mem[330] = 8'h00;
mem[331] = 8'h00;
mem[332] = 8'h00;
mem[333] = 8'h00;
mem[334] = 8'h00;
mem[335] = 8'h00;
mem[336] = 8'h00;
mem[337] = 8'h00;
mem[338] = 8'h00;
mem[339] = 8'h00;
mem[340] = 8'h00;
mem[341] = 8'h00;
mem[342] = 8'h00;
mem[343] = 8'h00;
mem[344] = 8'h00;
mem[345] = 8'h00;
mem[346] = 8'h00;
mem[347] = 8'h00;
mem[348] = 8'h00;
mem[349] = 8'h00;
mem[350] = 8'h00;
mem[351] = 8'h00;
mem[352] = 8'h00;
mem[353] = 8'h00;
mem[354] = 8'h00;
mem[355] = 8'h00;
mem[356] = 8'h00;
mem[357] = 8'h00;
mem[358] = 8'h00;
mem[359] = 8'h00;
mem[360] = 8'h00;
mem[361] = 8'h00;
mem[362] = 8'h00;
mem[363] = 8'h00;
mem[364] = 8'h00;
mem[365] = 8'h00;
mem[366] = 8'h00;
mem[367] = 8'h00;
mem[368] = 8'h00;
mem[369] = 8'h00;
mem[370] = 8'h00;
mem[371] = 8'h00;
mem[372] = 8'h00;
mem[373] = 8'h00;
mem[374] = 8'h00;
mem[375] = 8'h00;
mem[376] = 8'h00;
mem[377] = 8'h00;
mem[378] = 8'h00;
mem[379] = 8'h00;
mem[380] = 8'h00;
mem[381] = 8'h00;
mem[382] = 8'h00;
mem[383] = 8'h00;
mem[384] = 8'h00;
mem[385] = 8'h00;
mem[386] = 8'h00;
mem[387] = 8'h00;
mem[388] = 8'h00;
mem[389] = 8'h00;
mem[390] = 8'h00;
mem[391] = 8'h00;
mem[392] = 8'h00;
mem[393] = 8'h00;
mem[394] = 8'h00;
mem[395] = 8'h00;
mem[396] = 8'h00;
mem[397] = 8'h00;
mem[398] = 8'h00;
mem[399] = 8'h00;
mem[400] = 8'h00;
mem[401] = 8'h00;
mem[402] = 8'h00;
mem[403] = 8'h00;
mem[404] = 8'h00;
mem[405] = 8'h00;
mem[406] = 8'h00;
mem[407] = 8'h00;
mem[408] = 8'h00;
mem[409] = 8'h00;
mem[410] = 8'h00;
mem[411] = 8'h00;
mem[412] = 8'h00;
mem[413] = 8'h00;
mem[414] = 8'h00;
mem[415] = 8'h00;
mem[416] = 8'h00;
mem[417] = 8'h00;
mem[418] = 8'h00;
mem[419] = 8'h00;
mem[420] = 8'h00;
mem[421] = 8'h00;
mem[422] = 8'h00;
mem[423] = 8'h00;
mem[424] = 8'h00;
mem[425] = 8'h00;
mem[426] = 8'h00;
mem[427] = 8'h00;
mem[428] = 8'h00;
mem[429] = 8'h00;
mem[430] = 8'h00;
mem[431] = 8'h00;
mem[432] = 8'h00;
mem[433] = 8'h00;
mem[434] = 8'h00;
mem[435] = 8'h00;
mem[436] = 8'h00;
mem[437] = 8'h00;
mem[438] = 8'h00;
mem[439] = 8'h00;
mem[440] = 8'h00;
mem[441] = 8'h00;
mem[442] = 8'h00;
mem[443] = 8'h00;
mem[444] = 8'h00;
mem[445] = 8'h00;
mem[446] = 8'h00;
mem[447] = 8'h00;
mem[448] = 8'h00;
mem[449] = 8'h00;
mem[450] = 8'h00;
mem[451] = 8'h00;
mem[452] = 8'h00;
mem[453] = 8'h00;
mem[454] = 8'h00;
mem[455] = 8'h00;
mem[456] = 8'h00;
mem[457] = 8'h00;
mem[458] = 8'h00;
mem[459] = 8'h00;
mem[460] = 8'h00;
mem[461] = 8'h00;
mem[462] = 8'h00;
mem[463] = 8'h00;
mem[464] = 8'h00;
mem[465] = 8'h00;
mem[466] = 8'h00;
mem[467] = 8'h00;
mem[468] = 8'h00;
mem[469] = 8'h00;
mem[470] = 8'h00;
mem[471] = 8'h00;
mem[472] = 8'h00;
mem[473] = 8'h00;
mem[474] = 8'h00;
mem[475] = 8'h00;
mem[476] = 8'h00;
mem[477] = 8'h00;
mem[478] = 8'h00;
mem[479] = 8'h00;
mem[480] = 8'h00;
mem[481] = 8'h00;
mem[482] = 8'h00;
mem[483] = 8'h00;
mem[484] = 8'h00;
mem[485] = 8'h00;
mem[486] = 8'h00;
mem[487] = 8'h00;
mem[488] = 8'h00;
mem[489] = 8'h00;
mem[490] = 8'h00;
mem[491] = 8'h00;
mem[492] = 8'h00;
mem[493] = 8'h00;
mem[494] = 8'h00;
mem[495] = 8'h00;
mem[496] = 8'h00;
mem[497] = 8'h00;
mem[498] = 8'h00;
mem[499] = 8'h00;
mem[500] = 8'h00;
mem[501] = 8'h00;
mem[502] = 8'h00;
mem[503] = 8'h00;
mem[504] = 8'h00;
mem[505] = 8'h00;
mem[506] = 8'h00;
mem[507] = 8'h00;
mem[508] = 8'h00;
mem[509] = 8'h00;
mem[510] = 8'h00;
mem[511] = 8'h00;
mem[512] = 8'h00;
mem[513] = 8'h00;
mem[514] = 8'h00;
mem[515] = 8'h00;
mem[516] = 8'h00;
mem[517] = 8'h00;
mem[518] = 8'h00;
mem[519] = 8'h00;
mem[520] = 8'h00;
mem[521] = 8'h00;
mem[522] = 8'h00;
mem[523] = 8'h00;
mem[524] = 8'h00;
mem[525] = 8'h00;
mem[526] = 8'h00;
mem[527] = 8'h00;
mem[528] = 8'h00;
mem[529] = 8'h00;
mem[530] = 8'h00;
mem[531] = 8'h00;
mem[532] = 8'h00;
mem[533] = 8'h00;
mem[534] = 8'h00;
mem[535] = 8'h00;
mem[536] = 8'h00;
mem[537] = 8'h00;
mem[538] = 8'h00;
mem[539] = 8'h00;
mem[540] = 8'h00;
mem[541] = 8'h00;
mem[542] = 8'h00;
mem[543] = 8'h00;
mem[544] = 8'h00;
mem[545] = 8'h00;
mem[546] = 8'h00;
mem[547] = 8'h00;
mem[548] = 8'h00;
mem[549] = 8'h00;
mem[550] = 8'h00;
mem[551] = 8'h00;
mem[552] = 8'h00;
mem[553] = 8'h00;
mem[554] = 8'h00;
mem[555] = 8'h00;
mem[556] = 8'h00;
mem[557] = 8'h00;
mem[558] = 8'h00;
mem[559] = 8'h00;
mem[560] = 8'h00;
mem[561] = 8'h00;
mem[562] = 8'h00;
mem[563] = 8'h00;
mem[564] = 8'h00;
mem[565] = 8'h00;
mem[566] = 8'h00;
mem[567] = 8'h00;
mem[568] = 8'h00;
mem[569] = 8'h00;
mem[570] = 8'h00;
mem[571] = 8'h00;
mem[572] = 8'h00;
mem[573] = 8'h00;
mem[574] = 8'h00;
mem[575] = 8'h00;
mem[576] = 8'h00;
mem[577] = 8'h00;
mem[578] = 8'h00;
mem[579] = 8'h00;
mem[580] = 8'h00;
mem[581] = 8'h00;
mem[582] = 8'h00;
mem[583] = 8'h00;
mem[584] = 8'h00;
mem[585] = 8'h00;
mem[586] = 8'h00;
mem[587] = 8'h00;
mem[588] = 8'h00;
mem[589] = 8'h00;
mem[590] = 8'h00;
mem[591] = 8'h00;
mem[592] = 8'h00;
mem[593] = 8'h00;
mem[594] = 8'h00;
mem[595] = 8'h00;
mem[596] = 8'h00;
mem[597] = 8'h00;
mem[598] = 8'h00;
mem[599] = 8'h00;
mem[600] = 8'h00;
mem[601] = 8'h00;
mem[602] = 8'h00;
mem[603] = 8'h00;
mem[604] = 8'h00;
mem[605] = 8'h00;
mem[606] = 8'h00;
mem[607] = 8'h00;
mem[608] = 8'h00;
mem[609] = 8'h00;
mem[610] = 8'h00;
mem[611] = 8'h00;
mem[612] = 8'h00;
mem[613] = 8'h00;
mem[614] = 8'h00;
mem[615] = 8'h00;
mem[616] = 8'h00;
mem[617] = 8'h00;
mem[618] = 8'h00;
mem[619] = 8'h00;
mem[620] = 8'h00;
mem[621] = 8'h00;
mem[622] = 8'h00;
mem[623] = 8'h00;
mem[624] = 8'h00;
mem[625] = 8'h00;
mem[626] = 8'h00;
mem[627] = 8'h00;
mem[628] = 8'h00;
mem[629] = 8'h00;
mem[630] = 8'h00;
mem[631] = 8'h00;
mem[632] = 8'h00;
mem[633] = 8'h00;
mem[634] = 8'h00;
mem[635] = 8'h00;
mem[636] = 8'h00;
mem[637] = 8'h00;
mem[638] = 8'h00;
mem[639] = 8'h00;
mem[640] = 8'h00;
mem[641] = 8'h00;
mem[642] = 8'h00;
mem[643] = 8'h00;
mem[644] = 8'h00;
mem[645] = 8'h00;
mem[646] = 8'h00;
mem[647] = 8'h00;
mem[648] = 8'h00;
mem[649] = 8'h00;
mem[650] = 8'h00;
mem[651] = 8'h00;
mem[652] = 8'h00;
mem[653] = 8'h00;
mem[654] = 8'h00;
mem[655] = 8'h00;
mem[656] = 8'h00;
mem[657] = 8'h00;
mem[658] = 8'h00;
mem[659] = 8'h00;
mem[660] = 8'h00;
mem[661] = 8'h00;
mem[662] = 8'h00;
mem[663] = 8'h00;
mem[664] = 8'h00;
mem[665] = 8'h00;
mem[666] = 8'h00;
mem[667] = 8'h00;
mem[668] = 8'h00;
mem[669] = 8'h00;
mem[670] = 8'h00;
mem[671] = 8'h00;
mem[672] = 8'h00;
mem[673] = 8'h00;
mem[674] = 8'h00;
mem[675] = 8'h00;
mem[676] = 8'h00;
mem[677] = 8'h00;
mem[678] = 8'h00;
mem[679] = 8'h00;
mem[680] = 8'h00;
mem[681] = 8'h00;
mem[682] = 8'h00;
mem[683] = 8'h00;
mem[684] = 8'h00;
mem[685] = 8'h00;
mem[686] = 8'h00;
mem[687] = 8'h00;
mem[688] = 8'h00;
mem[689] = 8'h00;
mem[690] = 8'h00;
mem[691] = 8'h00;
mem[692] = 8'h00;
mem[693] = 8'h00;
mem[694] = 8'h00;
mem[695] = 8'h00;
mem[696] = 8'h00;
mem[697] = 8'h00;
mem[698] = 8'h00;
mem[699] = 8'h00;
mem[700] = 8'h00;
mem[701] = 8'h00;
mem[702] = 8'h00;
mem[703] = 8'h00;
mem[704] = 8'h00;
mem[705] = 8'h00;
mem[706] = 8'h00;
mem[707] = 8'h00;
mem[708] = 8'h00;
mem[709] = 8'h00;
mem[710] = 8'h00;
mem[711] = 8'h00;
mem[712] = 8'h00;
mem[713] = 8'h00;
mem[714] = 8'h00;
mem[715] = 8'h00;
mem[716] = 8'h00;
mem[717] = 8'h00;
mem[718] = 8'h00;
mem[719] = 8'h00;
mem[720] = 8'h00;
mem[721] = 8'h00;
mem[722] = 8'h00;
mem[723] = 8'h00;
mem[724] = 8'h00;
mem[725] = 8'h00;
mem[726] = 8'h00;
mem[727] = 8'h00;
mem[728] = 8'h00;
mem[729] = 8'h00;
mem[730] = 8'h00;
mem[731] = 8'h00;
mem[732] = 8'h00;
mem[733] = 8'h00;
mem[734] = 8'h00;
mem[735] = 8'h00;
mem[736] = 8'h00;
mem[737] = 8'h00;
mem[738] = 8'h00;
mem[739] = 8'h00;
mem[740] = 8'h00;
mem[741] = 8'h00;
mem[742] = 8'h00;
mem[743] = 8'h00;
mem[744] = 8'h00;
mem[745] = 8'h00;
mem[746] = 8'h00;
mem[747] = 8'h00;
mem[748] = 8'h00;
mem[749] = 8'h00;
mem[750] = 8'h00;
mem[751] = 8'h00;
mem[752] = 8'h00;
mem[753] = 8'h00;
mem[754] = 8'h00;
mem[755] = 8'h00;
mem[756] = 8'h00;
mem[757] = 8'h00;
mem[758] = 8'h00;
mem[759] = 8'h00;
mem[760] = 8'h00;
mem[761] = 8'h00;
mem[762] = 8'h00;
mem[763] = 8'h00;
mem[764] = 8'h00;
mem[765] = 8'h00;
mem[766] = 8'h00;
mem[767] = 8'h00;
mem[768] = 8'h00;
mem[769] = 8'h00;
mem[770] = 8'h00;
mem[771] = 8'h00;
mem[772] = 8'h00;
mem[773] = 8'h00;
mem[774] = 8'h00;
mem[775] = 8'h00;
mem[776] = 8'h00;
mem[777] = 8'h00;
mem[778] = 8'h00;
mem[779] = 8'h00;
mem[780] = 8'h00;
mem[781] = 8'h00;
mem[782] = 8'h00;
mem[783] = 8'h00;
mem[784] = 8'h00;
mem[785] = 8'h00;
mem[786] = 8'h00;
mem[787] = 8'h00;
mem[788] = 8'h00;
mem[789] = 8'h00;
mem[790] = 8'h00;
mem[791] = 8'h00;
mem[792] = 8'h00;
mem[793] = 8'h00;
mem[794] = 8'h00;
mem[795] = 8'h00;
mem[796] = 8'h00;
mem[797] = 8'h00;
mem[798] = 8'h00;
mem[799] = 8'h00;
mem[800] = 8'h00;
mem[801] = 8'h00;
mem[802] = 8'h00;
mem[803] = 8'h00;
mem[804] = 8'h00;
mem[805] = 8'h00;
mem[806] = 8'h00;
mem[807] = 8'h00;
mem[808] = 8'h00;
mem[809] = 8'h00;
mem[810] = 8'h00;
mem[811] = 8'h00;
mem[812] = 8'h00;
mem[813] = 8'h00;
mem[814] = 8'h00;
mem[815] = 8'h00;
mem[816] = 8'h00;
mem[817] = 8'h00;
mem[818] = 8'h00;
mem[819] = 8'h00;
mem[820] = 8'h00;
mem[821] = 8'h00;
mem[822] = 8'h00;
mem[823] = 8'h00;
mem[824] = 8'h00;
mem[825] = 8'h00;
mem[826] = 8'h00;
mem[827] = 8'h00;
mem[828] = 8'h00;
mem[829] = 8'h00;
mem[830] = 8'h00;
mem[831] = 8'h00;
mem[832] = 8'h00;
mem[833] = 8'h00;
mem[834] = 8'h00;
mem[835] = 8'h00;
mem[836] = 8'h00;
mem[837] = 8'h00;
mem[838] = 8'h00;
mem[839] = 8'h00;
mem[840] = 8'h00;
mem[841] = 8'h00;
mem[842] = 8'h00;
mem[843] = 8'h00;
mem[844] = 8'h00;
mem[845] = 8'h00;
mem[846] = 8'h00;
mem[847] = 8'h00;
mem[848] = 8'h00;
mem[849] = 8'h00;
mem[850] = 8'h00;
mem[851] = 8'h00;
mem[852] = 8'h00;
mem[853] = 8'h00;
mem[854] = 8'h00;
mem[855] = 8'h00;
mem[856] = 8'h00;
mem[857] = 8'h00;
mem[858] = 8'h00;
mem[859] = 8'h00;
mem[860] = 8'h00;
mem[861] = 8'h00;
mem[862] = 8'h00;
mem[863] = 8'h00;
mem[864] = 8'h00;
mem[865] = 8'h00;
mem[866] = 8'h00;
mem[867] = 8'h00;
mem[868] = 8'h00;
mem[869] = 8'h00;
mem[870] = 8'h00;
mem[871] = 8'h00;
mem[872] = 8'h00;
mem[873] = 8'h00;
mem[874] = 8'h00;
mem[875] = 8'h00;
mem[876] = 8'h00;
mem[877] = 8'h00;
mem[878] = 8'h00;
mem[879] = 8'h00;
mem[880] = 8'h00;
mem[881] = 8'h00;
mem[882] = 8'h00;
mem[883] = 8'h00;
mem[884] = 8'h00;
mem[885] = 8'h00;
mem[886] = 8'h00;
mem[887] = 8'h00;
mem[888] = 8'h00;
mem[889] = 8'h00;
mem[890] = 8'h00;
mem[891] = 8'h00;
mem[892] = 8'h00;
mem[893] = 8'h00;
mem[894] = 8'h00;
mem[895] = 8'h00;
mem[896] = 8'h00;
mem[897] = 8'h00;
mem[898] = 8'h00;
mem[899] = 8'h00;
mem[900] = 8'h00;
mem[901] = 8'h00;
mem[902] = 8'h00;
mem[903] = 8'h00;
mem[904] = 8'h00;
mem[905] = 8'h00;
mem[906] = 8'h00;
mem[907] = 8'h00;
mem[908] = 8'h00;
mem[909] = 8'h00;
mem[910] = 8'h00;
mem[911] = 8'h00;
mem[912] = 8'h00;
mem[913] = 8'h00;
mem[914] = 8'h00;
mem[915] = 8'h00;
mem[916] = 8'h00;
mem[917] = 8'h00;
mem[918] = 8'h00;
mem[919] = 8'h00;
mem[920] = 8'h00;
mem[921] = 8'h00;
mem[922] = 8'h00;
mem[923] = 8'h00;
mem[924] = 8'h00;
mem[925] = 8'h00;
mem[926] = 8'h00;
mem[927] = 8'h00;
mem[928] = 8'h00;
mem[929] = 8'h00;
mem[930] = 8'h00;
mem[931] = 8'h00;
mem[932] = 8'h00;
mem[933] = 8'h00;
mem[934] = 8'h00;
mem[935] = 8'h00;
mem[936] = 8'h00;
mem[937] = 8'h00;
mem[938] = 8'h00;
mem[939] = 8'h00;
mem[940] = 8'h00;
mem[941] = 8'h00;
mem[942] = 8'h00;
mem[943] = 8'h00;
mem[944] = 8'h00;
mem[945] = 8'h00;
mem[946] = 8'h00;
mem[947] = 8'h00;
mem[948] = 8'h00;
mem[949] = 8'h00;
mem[950] = 8'h00;
mem[951] = 8'h00;
mem[952] = 8'h00;
mem[953] = 8'h00;
mem[954] = 8'h00;
mem[955] = 8'h00;
mem[956] = 8'h00;
mem[957] = 8'h00;
mem[958] = 8'h00;
mem[959] = 8'h00;
mem[960] = 8'h00;
mem[961] = 8'h00;
mem[962] = 8'h00;
mem[963] = 8'h00;
mem[964] = 8'h00;
mem[965] = 8'h00;
mem[966] = 8'h00;
mem[967] = 8'h00;
mem[968] = 8'h00;
mem[969] = 8'h00;
mem[970] = 8'h00;
mem[971] = 8'h00;
mem[972] = 8'h00;
mem[973] = 8'h00;
mem[974] = 8'h00;
mem[975] = 8'h00;
mem[976] = 8'h00;
mem[977] = 8'h00;
mem[978] = 8'h00;
mem[979] = 8'h00;
mem[980] = 8'h00;
mem[981] = 8'h00;
mem[982] = 8'h00;
mem[983] = 8'h00;
mem[984] = 8'h00;
mem[985] = 8'h00;
mem[986] = 8'h00;
mem[987] = 8'h00;
mem[988] = 8'h00;
mem[989] = 8'h00;
mem[990] = 8'h00;
mem[991] = 8'h00;
mem[992] = 8'h00;
mem[993] = 8'h00;
mem[994] = 8'h00;
mem[995] = 8'h00;
mem[996] = 8'h00;
mem[997] = 8'h00;
mem[998] = 8'h00;
mem[999] = 8'h00;
mem[1000] = 8'h00;
mem[1001] = 8'h00;
mem[1002] = 8'h00;
mem[1003] = 8'h00;
mem[1004] = 8'h00;
mem[1005] = 8'h00;
mem[1006] = 8'h00;
mem[1007] = 8'h00;
mem[1008] = 8'h00;
mem[1009] = 8'h00;
mem[1010] = 8'h00;
mem[1011] = 8'h00;
mem[1012] = 8'h00;
mem[1013] = 8'h00;
mem[1014] = 8'h00;
mem[1015] = 8'h00;
mem[1016] = 8'h00;
mem[1017] = 8'h00;
mem[1018] = 8'h00;
mem[1019] = 8'h00;
mem[1020] = 8'h00;
mem[1021] = 8'h00;
mem[1022] = 8'h00;
mem[1023] = 8'h00;
mem[1024] = 8'hf0;
mem[1025] = 8'h01;
mem[1026] = 8'h02;
mem[1027] = 8'h03;
mem[1028] = 8'h04;
mem[1029] = 8'h05;
mem[1030] = 8'h06;
mem[1031] = 8'h07;
mem[1032] = 8'h08;
mem[1033] = 8'h09;
mem[1034] = 8'h0a;
mem[1035] = 8'h0b;
mem[1036] = 8'h0c;
mem[1037] = 8'h0d;
mem[1038] = 8'h0e;
mem[1039] = 8'h0f;
mem[1040] = 8'h0f;
mem[1041] = 8'h0e;
mem[1042] = 8'h0d;
mem[1043] = 8'h0c;
mem[1044] = 8'h0b;
mem[1045] = 8'h0a;
mem[1046] = 8'h09;
mem[1047] = 8'h08;
mem[1048] = 8'h07;
mem[1049] = 8'h06;
mem[1050] = 8'h05;
mem[1051] = 8'h04;
mem[1052] = 8'h03;
mem[1053] = 8'h02;
mem[1054] = 8'h01;
mem[1055] = 8'hf0;
mem[1056] = 8'h0f;
mem[1057] = 8'h0f;
mem[1058] = 8'h0f;
mem[1059] = 8'h0f;
mem[1060] = 8'h0f;
mem[1061] = 8'h0f;
mem[1062] = 8'h0f;
mem[1063] = 8'h0f;
mem[1064] = 8'h0f;
mem[1065] = 8'h0f;
mem[1066] = 8'h0f;
mem[1067] = 8'h0f;
mem[1068] = 8'h0f;
mem[1069] = 8'h0f;
mem[1070] = 8'h0f;
mem[1071] = 8'h0f;
mem[1072] = 8'h0f;
mem[1073] = 8'h0f;
mem[1074] = 8'h0f;
mem[1075] = 8'h0f;
mem[1076] = 8'h0f;
mem[1077] = 8'h0f;
mem[1078] = 8'h0f;
mem[1079] = 8'h0f;
mem[1080] = 8'h0f;
mem[1081] = 8'h0f;
mem[1082] = 8'h0f;
mem[1083] = 8'h0f;
mem[1084] = 8'h0f;
mem[1085] = 8'h0f;
mem[1086] = 8'h0f;
mem[1087] = 8'h0f;
mem[1088] = 8'h0f;
mem[1089] = 8'h0f;
mem[1090] = 8'h0f;
mem[1091] = 8'h0f;
mem[1092] = 8'h0f;
mem[1093] = 8'h0f;
mem[1094] = 8'h0f;
mem[1095] = 8'h0f;
mem[1096] = 8'h0f;
mem[1097] = 8'h0f;
mem[1098] = 8'h0f;
mem[1099] = 8'h0f;
mem[1100] = 8'h0f;
mem[1101] = 8'h0f;
mem[1102] = 8'h0f;
mem[1103] = 8'h0f;
mem[1104] = 8'h0f;
mem[1105] = 8'h0f;
mem[1106] = 8'h0f;
mem[1107] = 8'h0f;
mem[1108] = 8'h0f;
mem[1109] = 8'h0f;
mem[1110] = 8'h0f;
mem[1111] = 8'h0f;
mem[1112] = 8'h0f;
mem[1113] = 8'h0f;
mem[1114] = 8'h0f;
mem[1115] = 8'h0f;
mem[1116] = 8'h0f;
mem[1117] = 8'h0f;
mem[1118] = 8'h0f;
mem[1119] = 8'h0f;
mem[1120] = 8'h0f;
mem[1121] = 8'h0f;
mem[1122] = 8'h0f;
mem[1123] = 8'h0f;
mem[1124] = 8'h0f;
mem[1125] = 8'h0f;
mem[1126] = 8'h0f;
mem[1127] = 8'h0f;
mem[1128] = 8'h0f;
mem[1129] = 8'h0f;
mem[1130] = 8'h0f;
mem[1131] = 8'h0f;
mem[1132] = 8'h0f;
mem[1133] = 8'h0f;
mem[1134] = 8'h0f;
mem[1135] = 8'h0f;
mem[1136] = 8'h0f;
mem[1137] = 8'h0f;
mem[1138] = 8'h0f;
mem[1139] = 8'h0f;
mem[1140] = 8'h0f;
mem[1141] = 8'h0f;
mem[1142] = 8'h0f;
mem[1143] = 8'h0f;
mem[1144] = 8'h0f;
mem[1145] = 8'h0f;
mem[1146] = 8'h0f;
mem[1147] = 8'h0f;
mem[1148] = 8'h0f;
mem[1149] = 8'h0f;
mem[1150] = 8'h0f;
mem[1151] = 8'h0f;
mem[1152] = 8'h0f;
mem[1153] = 8'h0f;
mem[1154] = 8'h0f;
mem[1155] = 8'h0f;
mem[1156] = 8'h0f;
mem[1157] = 8'h0f;
mem[1158] = 8'h0f;
mem[1159] = 8'h0f;
mem[1160] = 8'h0f;
mem[1161] = 8'h0f;
mem[1162] = 8'h0f;
mem[1163] = 8'h0f;
mem[1164] = 8'h0f;
mem[1165] = 8'h0f;
mem[1166] = 8'h0f;
mem[1167] = 8'h0f;
mem[1168] = 8'h0f;
mem[1169] = 8'h0f;
mem[1170] = 8'h0f;
mem[1171] = 8'h0f;
mem[1172] = 8'h0f;
mem[1173] = 8'h0f;
mem[1174] = 8'h0f;
mem[1175] = 8'h0f;
mem[1176] = 8'h0f;
mem[1177] = 8'h0f;
mem[1178] = 8'h0f;
mem[1179] = 8'h0f;
mem[1180] = 8'h0f;
mem[1181] = 8'h0f;
mem[1182] = 8'h0f;
mem[1183] = 8'h0f;
mem[1184] = 8'h0f;
mem[1185] = 8'h0f;
mem[1186] = 8'h0f;
mem[1187] = 8'h0f;
mem[1188] = 8'h0f;
mem[1189] = 8'h0f;
mem[1190] = 8'h0f;
mem[1191] = 8'h0f;
mem[1192] = 8'h0f;
mem[1193] = 8'h0f;
mem[1194] = 8'h0f;
mem[1195] = 8'h0f;
mem[1196] = 8'h0f;
mem[1197] = 8'h0f;
mem[1198] = 8'h0f;
mem[1199] = 8'h0f;
mem[1200] = 8'h0f;
mem[1201] = 8'h0f;
mem[1202] = 8'h0f;
mem[1203] = 8'h0f;
mem[1204] = 8'h0f;
mem[1205] = 8'h0f;
mem[1206] = 8'h0f;
mem[1207] = 8'h0f;
mem[1208] = 8'h0f;
mem[1209] = 8'h0f;
mem[1210] = 8'h0f;
mem[1211] = 8'h0f;
mem[1212] = 8'h0f;
mem[1213] = 8'h0f;
mem[1214] = 8'h0f;
mem[1215] = 8'h0f;
mem[1216] = 8'h0f;
mem[1217] = 8'h0f;
mem[1218] = 8'h0f;
mem[1219] = 8'h0f;
mem[1220] = 8'h0f;
mem[1221] = 8'h0f;
mem[1222] = 8'h0f;
mem[1223] = 8'h0f;
mem[1224] = 8'h0f;
mem[1225] = 8'h0f;
mem[1226] = 8'h0f;
mem[1227] = 8'h0f;
mem[1228] = 8'h0f;
mem[1229] = 8'h0f;
mem[1230] = 8'h0f;
mem[1231] = 8'h0f;
mem[1232] = 8'h0f;
mem[1233] = 8'h0f;
mem[1234] = 8'h0f;
mem[1235] = 8'h0f;
mem[1236] = 8'h0f;
mem[1237] = 8'h0f;
mem[1238] = 8'h0f;
mem[1239] = 8'h0f;
mem[1240] = 8'h0f;
mem[1241] = 8'h0f;
mem[1242] = 8'h0f;
mem[1243] = 8'h0f;
mem[1244] = 8'h0f;
mem[1245] = 8'h0f;
mem[1246] = 8'h0f;
mem[1247] = 8'h0f;
mem[1248] = 8'h0f;
mem[1249] = 8'h0f;
mem[1250] = 8'h0f;
mem[1251] = 8'h0f;
mem[1252] = 8'h0f;
mem[1253] = 8'h0f;
mem[1254] = 8'h0f;
mem[1255] = 8'h0f;
mem[1256] = 8'h0f;
mem[1257] = 8'h0f;
mem[1258] = 8'h0f;
mem[1259] = 8'h0f;
mem[1260] = 8'h0f;
mem[1261] = 8'h0f;
mem[1262] = 8'h0f;
mem[1263] = 8'h0f;
mem[1264] = 8'h0f;
mem[1265] = 8'h0f;
mem[1266] = 8'h0f;
mem[1267] = 8'h0f;
mem[1268] = 8'h0f;
mem[1269] = 8'h0f;
mem[1270] = 8'h0f;
mem[1271] = 8'h0f;
mem[1272] = 8'h0f;
mem[1273] = 8'h0f;
mem[1274] = 8'h0f;
mem[1275] = 8'h0f;
mem[1276] = 8'h0f;
mem[1277] = 8'h0f;
mem[1278] = 8'h0f;
mem[1279] = 8'h0f;
mem[1280] = 8'h0f;
mem[1281] = 8'h0f;
mem[1282] = 8'h0f;
mem[1283] = 8'h0f;
mem[1284] = 8'h0f;
mem[1285] = 8'h0f;
mem[1286] = 8'h0f;
mem[1287] = 8'h0f;
mem[1288] = 8'h0f;
mem[1289] = 8'h0f;
mem[1290] = 8'h0f;
mem[1291] = 8'h0f;
mem[1292] = 8'h0f;
mem[1293] = 8'h0f;
mem[1294] = 8'h0f;
mem[1295] = 8'h0f;
mem[1296] = 8'h0f;
mem[1297] = 8'h0f;
mem[1298] = 8'h0f;
mem[1299] = 8'h0f;
mem[1300] = 8'h0f;
mem[1301] = 8'h0f;
mem[1302] = 8'h0f;
mem[1303] = 8'h0f;
mem[1304] = 8'h0f;
mem[1305] = 8'h0f;
mem[1306] = 8'h0f;
mem[1307] = 8'h0f;
mem[1308] = 8'h0f;
mem[1309] = 8'h0f;
mem[1310] = 8'h0f;
mem[1311] = 8'h0f;
mem[1312] = 8'h0f;
mem[1313] = 8'h0f;
mem[1314] = 8'h0f;
mem[1315] = 8'h0f;
mem[1316] = 8'h0f;
mem[1317] = 8'h0f;
mem[1318] = 8'h0f;
mem[1319] = 8'h0f;
mem[1320] = 8'h0f;
mem[1321] = 8'h0f;
mem[1322] = 8'h0f;
mem[1323] = 8'h0f;
mem[1324] = 8'h0f;
mem[1325] = 8'h0f;
mem[1326] = 8'h0f;
mem[1327] = 8'h0f;
mem[1328] = 8'h0f;
mem[1329] = 8'h0f;
mem[1330] = 8'h0f;
mem[1331] = 8'h0f;
mem[1332] = 8'h0f;
mem[1333] = 8'h0f;
mem[1334] = 8'h0f;
mem[1335] = 8'h0f;
mem[1336] = 8'h0f;
mem[1337] = 8'h0f;
mem[1338] = 8'h0f;
mem[1339] = 8'h0f;
mem[1340] = 8'h0f;
mem[1341] = 8'h0f;
mem[1342] = 8'h0f;
mem[1343] = 8'h0f;
mem[1344] = 8'h0f;
mem[1345] = 8'h0f;
mem[1346] = 8'h0f;
mem[1347] = 8'h0f;
mem[1348] = 8'h0f;
mem[1349] = 8'h0f;
mem[1350] = 8'h0f;
mem[1351] = 8'h0f;
mem[1352] = 8'h0f;
mem[1353] = 8'h0f;
mem[1354] = 8'h0f;
mem[1355] = 8'h0f;
mem[1356] = 8'h0f;
mem[1357] = 8'h0f;
mem[1358] = 8'h0f;
mem[1359] = 8'h0f;
mem[1360] = 8'h0f;
mem[1361] = 8'h0f;
mem[1362] = 8'h0f;
mem[1363] = 8'h0f;
mem[1364] = 8'h0f;
mem[1365] = 8'h0f;
mem[1366] = 8'h0f;
mem[1367] = 8'h0f;
mem[1368] = 8'h0f;
mem[1369] = 8'h0f;
mem[1370] = 8'h0f;
mem[1371] = 8'h0f;
mem[1372] = 8'h0f;
mem[1373] = 8'h0f;
mem[1374] = 8'h0f;
mem[1375] = 8'h0f;
mem[1376] = 8'h0f;
mem[1377] = 8'h0f;
mem[1378] = 8'h0f;
mem[1379] = 8'h0f;
mem[1380] = 8'h0f;
mem[1381] = 8'h0f;
mem[1382] = 8'h0f;
mem[1383] = 8'h0f;
mem[1384] = 8'h0f;
mem[1385] = 8'h0f;
mem[1386] = 8'h0f;
mem[1387] = 8'h0f;
mem[1388] = 8'h0f;
mem[1389] = 8'h0f;
mem[1390] = 8'h0f;
mem[1391] = 8'h0f;
mem[1392] = 8'h0f;
mem[1393] = 8'h0f;
mem[1394] = 8'h0f;
mem[1395] = 8'h0f;
mem[1396] = 8'h0f;
mem[1397] = 8'h0f;
mem[1398] = 8'h0f;
mem[1399] = 8'h0f;
mem[1400] = 8'h0f;
mem[1401] = 8'h0f;
mem[1402] = 8'h0f;
mem[1403] = 8'h0f;
mem[1404] = 8'h0f;
mem[1405] = 8'h0f;
mem[1406] = 8'h0f;
mem[1407] = 8'h0f;
mem[1408] = 8'h0f;
mem[1409] = 8'h0f;
mem[1410] = 8'h0f;
mem[1411] = 8'h0f;
mem[1412] = 8'h0f;
mem[1413] = 8'h0f;
mem[1414] = 8'h0f;
mem[1415] = 8'h0f;
mem[1416] = 8'h0f;
mem[1417] = 8'h0f;
mem[1418] = 8'h0f;
mem[1419] = 8'h0f;
mem[1420] = 8'h0f;
mem[1421] = 8'h0f;
mem[1422] = 8'h0f;
mem[1423] = 8'h0f;
mem[1424] = 8'h0f;
mem[1425] = 8'h0f;
mem[1426] = 8'h0f;
mem[1427] = 8'h0f;
mem[1428] = 8'h0f;
mem[1429] = 8'h0f;
mem[1430] = 8'h0f;
mem[1431] = 8'h0f;
mem[1432] = 8'h0f;
mem[1433] = 8'h0f;
mem[1434] = 8'h0f;
mem[1435] = 8'h0f;
mem[1436] = 8'h0f;
mem[1437] = 8'h0f;
mem[1438] = 8'h0f;
mem[1439] = 8'h0f;
mem[1440] = 8'h0f;
mem[1441] = 8'h0f;
mem[1442] = 8'h0f;
mem[1443] = 8'h0f;
mem[1444] = 8'h0f;
mem[1445] = 8'h0f;
mem[1446] = 8'h0f;
mem[1447] = 8'h0f;
mem[1448] = 8'h0f;
mem[1449] = 8'h0f;
mem[1450] = 8'h0f;
mem[1451] = 8'h0f;
mem[1452] = 8'h0f;
mem[1453] = 8'h0f;
mem[1454] = 8'h0f;
mem[1455] = 8'h0f;
mem[1456] = 8'h0f;
mem[1457] = 8'h0f;
mem[1458] = 8'h0f;
mem[1459] = 8'h0f;
mem[1460] = 8'h0f;
mem[1461] = 8'h0f;
mem[1462] = 8'h0f;
mem[1463] = 8'h0f;
mem[1464] = 8'h0f;
mem[1465] = 8'h0f;
mem[1466] = 8'h0f;
mem[1467] = 8'h0f;
mem[1468] = 8'h0f;
mem[1469] = 8'h0f;
mem[1470] = 8'h0f;
mem[1471] = 8'h0f;
mem[1472] = 8'h0f;
mem[1473] = 8'h0f;
mem[1474] = 8'h0f;
mem[1475] = 8'h0f;
mem[1476] = 8'h0f;
mem[1477] = 8'h0f;
mem[1478] = 8'h0f;
mem[1479] = 8'h0f;
mem[1480] = 8'h0f;
mem[1481] = 8'h0f;
mem[1482] = 8'h0f;
mem[1483] = 8'h0f;
mem[1484] = 8'h0f;
mem[1485] = 8'h0f;
mem[1486] = 8'h0f;
mem[1487] = 8'h0f;
mem[1488] = 8'h0f;
mem[1489] = 8'h0f;
mem[1490] = 8'h0f;
mem[1491] = 8'h0f;
mem[1492] = 8'h0f;
mem[1493] = 8'h0f;
mem[1494] = 8'h0f;
mem[1495] = 8'h0f;
mem[1496] = 8'h0f;
mem[1497] = 8'h0f;
mem[1498] = 8'h0f;
mem[1499] = 8'h0f;
mem[1500] = 8'h0f;
mem[1501] = 8'h0f;
mem[1502] = 8'h0f;
mem[1503] = 8'h0f;
mem[1504] = 8'h0f;
mem[1505] = 8'h0f;
mem[1506] = 8'h0f;
mem[1507] = 8'h0f;
mem[1508] = 8'h0f;
mem[1509] = 8'h0f;
mem[1510] = 8'h0f;
mem[1511] = 8'h0f;
mem[1512] = 8'h0f;
mem[1513] = 8'h0f;
mem[1514] = 8'h0f;
mem[1515] = 8'h0f;
mem[1516] = 8'h0f;
mem[1517] = 8'h0f;
mem[1518] = 8'h0f;
mem[1519] = 8'h0f;
mem[1520] = 8'h0f;
mem[1521] = 8'h0f;
mem[1522] = 8'h0f;
mem[1523] = 8'h0f;
mem[1524] = 8'h0f;
mem[1525] = 8'h0f;
mem[1526] = 8'h0f;
mem[1527] = 8'h0f;
mem[1528] = 8'h0f;
mem[1529] = 8'h0f;
mem[1530] = 8'h0f;
mem[1531] = 8'h0f;
mem[1532] = 8'h0f;
mem[1533] = 8'h0f;
mem[1534] = 8'h0f;
mem[1535] = 8'h0f;
mem[1536] = 8'h0f;
mem[1537] = 8'h0f;
mem[1538] = 8'h0f;
mem[1539] = 8'h0f;
mem[1540] = 8'h0f;
mem[1541] = 8'h0f;
mem[1542] = 8'h0f;
mem[1543] = 8'h0f;
mem[1544] = 8'h0f;
mem[1545] = 8'h0f;
mem[1546] = 8'h0f;
mem[1547] = 8'h0f;
mem[1548] = 8'h0f;
mem[1549] = 8'h0f;
mem[1550] = 8'h0f;
mem[1551] = 8'h0f;
mem[1552] = 8'h0f;
mem[1553] = 8'h0f;
mem[1554] = 8'h0f;
mem[1555] = 8'h0f;
mem[1556] = 8'h0f;
mem[1557] = 8'h0f;
mem[1558] = 8'h0f;
mem[1559] = 8'h0f;
mem[1560] = 8'h0f;
mem[1561] = 8'h0f;
mem[1562] = 8'h0f;
mem[1563] = 8'h0f;
mem[1564] = 8'h0f;
mem[1565] = 8'h0f;
mem[1566] = 8'h0f;
mem[1567] = 8'h0f;
mem[1568] = 8'h0f;
mem[1569] = 8'h0f;
mem[1570] = 8'h0f;
mem[1571] = 8'h0f;
mem[1572] = 8'h0f;
mem[1573] = 8'h0f;
mem[1574] = 8'h0f;
mem[1575] = 8'h0f;
mem[1576] = 8'h0f;
mem[1577] = 8'h0f;
mem[1578] = 8'h0f;
mem[1579] = 8'h0f;
mem[1580] = 8'h0f;
mem[1581] = 8'h0f;
mem[1582] = 8'h0f;
mem[1583] = 8'h0f;
mem[1584] = 8'h0f;
mem[1585] = 8'h0f;
mem[1586] = 8'h0f;
mem[1587] = 8'h0f;
mem[1588] = 8'h0f;
mem[1589] = 8'h0f;
mem[1590] = 8'h0f;
mem[1591] = 8'h0f;
mem[1592] = 8'h0f;
mem[1593] = 8'h0f;
mem[1594] = 8'h0f;
mem[1595] = 8'h0f;
mem[1596] = 8'h0f;
mem[1597] = 8'h0f;
mem[1598] = 8'h0f;
mem[1599] = 8'h0f;
mem[1600] = 8'h0f;
mem[1601] = 8'h0f;
mem[1602] = 8'h0f;
mem[1603] = 8'h0f;
mem[1604] = 8'h0f;
mem[1605] = 8'h0f;
mem[1606] = 8'h0f;
mem[1607] = 8'h0f;
mem[1608] = 8'h0f;
mem[1609] = 8'h0f;
mem[1610] = 8'h0f;
mem[1611] = 8'h0f;
mem[1612] = 8'h0f;
mem[1613] = 8'h0f;
mem[1614] = 8'h0f;
mem[1615] = 8'h0f;
mem[1616] = 8'h0f;
mem[1617] = 8'h0f;
mem[1618] = 8'h0f;
mem[1619] = 8'h0f;
mem[1620] = 8'h0f;
mem[1621] = 8'h0f;
mem[1622] = 8'h0f;
mem[1623] = 8'h0f;
mem[1624] = 8'h0f;
mem[1625] = 8'h0f;
mem[1626] = 8'h0f;
mem[1627] = 8'h0f;
mem[1628] = 8'h0f;
mem[1629] = 8'h0f;
mem[1630] = 8'h0f;
mem[1631] = 8'h0f;
mem[1632] = 8'h0f;
mem[1633] = 8'h0f;
mem[1634] = 8'h0f;
mem[1635] = 8'h0f;
mem[1636] = 8'h0f;
mem[1637] = 8'h0f;
mem[1638] = 8'h0f;
mem[1639] = 8'h0f;
mem[1640] = 8'h0f;
mem[1641] = 8'h0f;
mem[1642] = 8'h0f;
mem[1643] = 8'h0f;
mem[1644] = 8'h0f;
mem[1645] = 8'h0f;
mem[1646] = 8'h0f;
mem[1647] = 8'h0f;
mem[1648] = 8'h0f;
mem[1649] = 8'h0f;
mem[1650] = 8'h0f;
mem[1651] = 8'h0f;
mem[1652] = 8'h0f;
mem[1653] = 8'h0f;
mem[1654] = 8'h0f;
mem[1655] = 8'h0f;
mem[1656] = 8'h0f;
mem[1657] = 8'h0f;
mem[1658] = 8'h0f;
mem[1659] = 8'h0f;
mem[1660] = 8'h0f;
mem[1661] = 8'h0f;
mem[1662] = 8'h0f;
mem[1663] = 8'h0f;
mem[1664] = 8'h0f;
mem[1665] = 8'h0f;
mem[1666] = 8'h0f;
mem[1667] = 8'h0f;
mem[1668] = 8'h0f;
mem[1669] = 8'h0f;
mem[1670] = 8'h0f;
mem[1671] = 8'h0f;
mem[1672] = 8'h0f;
mem[1673] = 8'h0f;
mem[1674] = 8'h0f;
mem[1675] = 8'h0f;
mem[1676] = 8'h0f;
mem[1677] = 8'h0f;
mem[1678] = 8'h0f;
mem[1679] = 8'h0f;
mem[1680] = 8'h0f;
mem[1681] = 8'h0f;
mem[1682] = 8'h0f;
mem[1683] = 8'h0f;
mem[1684] = 8'h0f;
mem[1685] = 8'h0f;
mem[1686] = 8'h0f;
mem[1687] = 8'h0f;
mem[1688] = 8'h0f;
mem[1689] = 8'h0f;
mem[1690] = 8'h0f;
mem[1691] = 8'h0f;
mem[1692] = 8'h0f;
mem[1693] = 8'h0f;
mem[1694] = 8'h0f;
mem[1695] = 8'h0f;
mem[1696] = 8'h0f;
mem[1697] = 8'h0f;
mem[1698] = 8'h0f;
mem[1699] = 8'h0f;
mem[1700] = 8'h0f;
mem[1701] = 8'h0f;
mem[1702] = 8'h0f;
mem[1703] = 8'h0f;
mem[1704] = 8'h0f;
mem[1705] = 8'h0f;
mem[1706] = 8'h0f;
mem[1707] = 8'h0f;
mem[1708] = 8'h0f;
mem[1709] = 8'h0f;
mem[1710] = 8'h0f;
mem[1711] = 8'h0f;
mem[1712] = 8'h0f;
mem[1713] = 8'h0f;
mem[1714] = 8'h0f;
mem[1715] = 8'h0f;
mem[1716] = 8'h0f;
mem[1717] = 8'h0f;
mem[1718] = 8'h0f;
mem[1719] = 8'h0f;
mem[1720] = 8'h0f;
mem[1721] = 8'h0f;
mem[1722] = 8'h0f;
mem[1723] = 8'h0f;
mem[1724] = 8'h0f;
mem[1725] = 8'h0f;
mem[1726] = 8'h0f;
mem[1727] = 8'h0f;
mem[1728] = 8'h0f;
mem[1729] = 8'h0f;
mem[1730] = 8'h0f;
mem[1731] = 8'h0f;
mem[1732] = 8'h0f;
mem[1733] = 8'h0f;
mem[1734] = 8'h0f;
mem[1735] = 8'h0f;
mem[1736] = 8'h0f;
mem[1737] = 8'h0f;
mem[1738] = 8'h0f;
mem[1739] = 8'h0f;
mem[1740] = 8'h0f;
mem[1741] = 8'h0f;
mem[1742] = 8'h0f;
mem[1743] = 8'h0f;
mem[1744] = 8'h0f;
mem[1745] = 8'h0f;
mem[1746] = 8'h0f;
mem[1747] = 8'h0f;
mem[1748] = 8'h0f;
mem[1749] = 8'h0f;
mem[1750] = 8'h0f;
mem[1751] = 8'h0f;
mem[1752] = 8'h0f;
mem[1753] = 8'h0f;
mem[1754] = 8'h0f;
mem[1755] = 8'h0f;
mem[1756] = 8'h0f;
mem[1757] = 8'h0f;
mem[1758] = 8'h0f;
mem[1759] = 8'h0f;
mem[1760] = 8'h0f;
mem[1761] = 8'h0f;
mem[1762] = 8'h0f;
mem[1763] = 8'h0f;
mem[1764] = 8'h0f;
mem[1765] = 8'h0f;
mem[1766] = 8'h0f;
mem[1767] = 8'h0f;
mem[1768] = 8'h0f;
mem[1769] = 8'h0f;
mem[1770] = 8'h0f;
mem[1771] = 8'h0f;
mem[1772] = 8'h0f;
mem[1773] = 8'h0f;
mem[1774] = 8'h0f;
mem[1775] = 8'h0f;
mem[1776] = 8'h0f;
mem[1777] = 8'h0f;
mem[1778] = 8'h0f;
mem[1779] = 8'h0f;
mem[1780] = 8'h0f;
mem[1781] = 8'h0f;
mem[1782] = 8'h0f;
mem[1783] = 8'h0f;
mem[1784] = 8'h0f;
mem[1785] = 8'h0f;
mem[1786] = 8'h0f;
mem[1787] = 8'h0f;
mem[1788] = 8'h0f;
mem[1789] = 8'h0f;
mem[1790] = 8'h0f;
mem[1791] = 8'h0f;
mem[1792] = 8'h0f;
mem[1793] = 8'h0f;
mem[1794] = 8'h0f;
mem[1795] = 8'h0f;
mem[1796] = 8'h0f;
mem[1797] = 8'h0f;
mem[1798] = 8'h0f;
mem[1799] = 8'h0f;
mem[1800] = 8'h0f;
mem[1801] = 8'h0f;
mem[1802] = 8'h0f;
mem[1803] = 8'h0f;
mem[1804] = 8'h0f;
mem[1805] = 8'h0f;
mem[1806] = 8'h0f;
mem[1807] = 8'h0f;
mem[1808] = 8'h0f;
mem[1809] = 8'h0f;
mem[1810] = 8'h0f;
mem[1811] = 8'h0f;
mem[1812] = 8'h0f;
mem[1813] = 8'h0f;
mem[1814] = 8'h0f;
mem[1815] = 8'h0f;
mem[1816] = 8'h0f;
mem[1817] = 8'h0f;
mem[1818] = 8'h0f;
mem[1819] = 8'h0f;
mem[1820] = 8'h0f;
mem[1821] = 8'h0f;
mem[1822] = 8'h0f;
mem[1823] = 8'h0f;
mem[1824] = 8'h0f;
mem[1825] = 8'h0f;
mem[1826] = 8'h0f;
mem[1827] = 8'h0f;
mem[1828] = 8'h0f;
mem[1829] = 8'h0f;
mem[1830] = 8'h0f;
mem[1831] = 8'h0f;
mem[1832] = 8'h0f;
mem[1833] = 8'h0f;
mem[1834] = 8'h0f;
mem[1835] = 8'h0f;
mem[1836] = 8'h0f;
mem[1837] = 8'h0f;
mem[1838] = 8'h0f;
mem[1839] = 8'h0f;
mem[1840] = 8'h0f;
mem[1841] = 8'h0f;
mem[1842] = 8'h0f;
mem[1843] = 8'h0f;
mem[1844] = 8'h0f;
mem[1845] = 8'h0f;
mem[1846] = 8'h0f;
mem[1847] = 8'h0f;
mem[1848] = 8'h0f;
mem[1849] = 8'h0f;
mem[1850] = 8'h0f;
mem[1851] = 8'h0f;
mem[1852] = 8'h0f;
mem[1853] = 8'h0f;
mem[1854] = 8'h0f;
mem[1855] = 8'h0f;
mem[1856] = 8'h0f;
mem[1857] = 8'h0f;
mem[1858] = 8'h0f;
mem[1859] = 8'h0f;
mem[1860] = 8'h0f;
mem[1861] = 8'h0f;
mem[1862] = 8'h0f;
mem[1863] = 8'h0f;
mem[1864] = 8'h0f;
mem[1865] = 8'h0f;
mem[1866] = 8'h0f;
mem[1867] = 8'h0f;
mem[1868] = 8'h0f;
mem[1869] = 8'h0f;
mem[1870] = 8'h0f;
mem[1871] = 8'h0f;
mem[1872] = 8'h0f;
mem[1873] = 8'h0f;
mem[1874] = 8'h0f;
mem[1875] = 8'h0f;
mem[1876] = 8'h0f;
mem[1877] = 8'h0f;
mem[1878] = 8'h0f;
mem[1879] = 8'h0f;
mem[1880] = 8'h0f;
mem[1881] = 8'h0f;
mem[1882] = 8'h0f;
mem[1883] = 8'h0f;
mem[1884] = 8'h0f;
mem[1885] = 8'h0f;
mem[1886] = 8'h0f;
mem[1887] = 8'h0f;
mem[1888] = 8'h0f;
mem[1889] = 8'h0f;
mem[1890] = 8'h0f;
mem[1891] = 8'h0f;
mem[1892] = 8'h0f;
mem[1893] = 8'h0f;
mem[1894] = 8'h0f;
mem[1895] = 8'h0f;
mem[1896] = 8'h0f;
mem[1897] = 8'h0f;
mem[1898] = 8'h0f;
mem[1899] = 8'h0f;
mem[1900] = 8'h0f;
mem[1901] = 8'h0f;
mem[1902] = 8'h0f;
mem[1903] = 8'h0f;
mem[1904] = 8'h0f;
mem[1905] = 8'h0f;
mem[1906] = 8'h0f;
mem[1907] = 8'h0f;
mem[1908] = 8'h0f;
mem[1909] = 8'h0f;
mem[1910] = 8'h0f;
mem[1911] = 8'h0f;
mem[1912] = 8'h0f;
mem[1913] = 8'h0f;
mem[1914] = 8'h0f;
mem[1915] = 8'h0f;
mem[1916] = 8'h0f;
mem[1917] = 8'h0f;
mem[1918] = 8'h0f;
mem[1919] = 8'h0f;
mem[1920] = 8'h0f;
mem[1921] = 8'h0f;
mem[1922] = 8'h0f;
mem[1923] = 8'h0f;
mem[1924] = 8'h0f;
mem[1925] = 8'h0f;
mem[1926] = 8'h0f;
mem[1927] = 8'h0f;
mem[1928] = 8'h0f;
mem[1929] = 8'h0f;
mem[1930] = 8'h0f;
mem[1931] = 8'h0f;
mem[1932] = 8'h0f;
mem[1933] = 8'h0f;
mem[1934] = 8'h0f;
mem[1935] = 8'h0f;
mem[1936] = 8'h0f;
mem[1937] = 8'h0f;
mem[1938] = 8'h0f;
mem[1939] = 8'h0f;
mem[1940] = 8'h0f;
mem[1941] = 8'h0f;
mem[1942] = 8'h0f;
mem[1943] = 8'h0f;
mem[1944] = 8'h0f;
mem[1945] = 8'h0f;
mem[1946] = 8'h0f;
mem[1947] = 8'h0f;
mem[1948] = 8'h0f;
mem[1949] = 8'h0f;
mem[1950] = 8'h0f;
mem[1951] = 8'h0f;
mem[1952] = 8'h0f;
mem[1953] = 8'h0f;
mem[1954] = 8'h0f;
mem[1955] = 8'h0f;
mem[1956] = 8'h0f;
mem[1957] = 8'h0f;
mem[1958] = 8'h0f;
mem[1959] = 8'h0f;
mem[1960] = 8'h0f;
mem[1961] = 8'h0f;
mem[1962] = 8'h0f;
mem[1963] = 8'h0f;
mem[1964] = 8'h0f;
mem[1965] = 8'h0f;
mem[1966] = 8'h0f;
mem[1967] = 8'h0f;
mem[1968] = 8'h0f;
mem[1969] = 8'h0f;
mem[1970] = 8'h0f;
mem[1971] = 8'h0f;
mem[1972] = 8'h0f;
mem[1973] = 8'h0f;
mem[1974] = 8'h0f;
mem[1975] = 8'h0f;
mem[1976] = 8'h0f;
mem[1977] = 8'h0f;
mem[1978] = 8'h0f;
mem[1979] = 8'h0f;
mem[1980] = 8'h0f;
mem[1981] = 8'h0f;
mem[1982] = 8'h0f;
mem[1983] = 8'h0f;
mem[1984] = 8'h0f;
mem[1985] = 8'h0f;
mem[1986] = 8'h0f;
mem[1987] = 8'h0f;
mem[1988] = 8'h0f;
mem[1989] = 8'h0f;
mem[1990] = 8'h0f;
mem[1991] = 8'h0f;
mem[1992] = 8'h0f;
mem[1993] = 8'h0f;
mem[1994] = 8'h0f;
mem[1995] = 8'h0f;
mem[1996] = 8'h0f;
mem[1997] = 8'h0f;
mem[1998] = 8'h0f;
mem[1999] = 8'h0f;
mem[2000] = 8'h0f;
mem[2001] = 8'h0f;
mem[2002] = 8'h0f;
mem[2003] = 8'h0f;
mem[2004] = 8'h0f;
mem[2005] = 8'h0f;
mem[2006] = 8'h0f;
mem[2007] = 8'h0f;
mem[2008] = 8'h0f;
mem[2009] = 8'h0f;
mem[2010] = 8'h0f;
mem[2011] = 8'h0f;
mem[2012] = 8'h0f;
mem[2013] = 8'h0f;
mem[2014] = 8'h0f;
mem[2015] = 8'h0f;
mem[2016] = 8'h0f;
mem[2017] = 8'h0f;
mem[2018] = 8'h0f;
mem[2019] = 8'h0f;
mem[2020] = 8'h0f;
mem[2021] = 8'h0f;
mem[2022] = 8'h0f;
mem[2023] = 8'h0f;
mem[2024] = 8'h0f;
mem[2025] = 8'h0f;
mem[2026] = 8'h0f;
mem[2027] = 8'h0f;
mem[2028] = 8'h0f;
mem[2029] = 8'h0f;
mem[2030] = 8'h0f;
mem[2031] = 8'h0f;
mem[2032] = 8'h0f;
mem[2033] = 8'h0f;
mem[2034] = 8'h0f;
mem[2035] = 8'h0f;
mem[2036] = 8'h0f;
mem[2037] = 8'h0f;
mem[2038] = 8'h0f;
mem[2039] = 8'h0f;
mem[2040] = 8'h0f;
mem[2041] = 8'h0f;
mem[2042] = 8'h0f;
mem[2043] = 8'h0f;
mem[2044] = 8'h0f;
mem[2045] = 8'h0f;
mem[2046] = 8'h0f;
mem[2047] = 8'h0f;
mem[2048] = 8'h00;
mem[2049] = 8'h00;
mem[2050] = 8'h00;
mem[2051] = 8'h00;
mem[2052] = 8'h00;
mem[2053] = 8'h00;
mem[2054] = 8'h00;
mem[2055] = 8'h00;
mem[2056] = 8'h01;
mem[2057] = 8'h03;
mem[2058] = 8'h03;
mem[2059] = 8'h06;
mem[2060] = 8'h06;
mem[2061] = 8'h0c;
mem[2062] = 8'h0c;
mem[2063] = 8'h18;
mem[2064] = 8'he0;
mem[2065] = 8'h38;
mem[2066] = 8'h0e;
mem[2067] = 8'h03;
mem[2068] = 8'h0e;
mem[2069] = 8'h38;
mem[2070] = 8'he0;
mem[2071] = 8'h00;
mem[2072] = 8'h07;
mem[2073] = 8'h1c;
mem[2074] = 8'h70;
mem[2075] = 8'hc0;
mem[2076] = 8'h30;
mem[2077] = 8'h1c;
mem[2078] = 8'h07;
mem[2079] = 8'h00;
mem[2080] = 8'hc3;
mem[2081] = 8'hc3;
mem[2082] = 8'h66;
mem[2083] = 8'h66;
mem[2084] = 8'h3c;
mem[2085] = 8'h3c;
mem[2086] = 8'h18;
mem[2087] = 8'h18;
mem[2088] = 8'h18;
mem[2089] = 8'h18;
mem[2090] = 8'h3c;
mem[2091] = 8'h3c;
mem[2092] = 8'h66;
mem[2093] = 8'h66;
mem[2094] = 8'hc3;
mem[2095] = 8'hc3;
mem[2096] = 8'h00;
mem[2097] = 8'h00;
mem[2098] = 8'h00;
mem[2099] = 8'h10;
mem[2100] = 8'h00;
mem[2101] = 8'h00;
mem[2102] = 8'h00;
mem[2103] = 8'h00;
mem[2104] = 8'h00;
mem[2105] = 8'h3f;
mem[2106] = 8'h3f;
mem[2107] = 8'h3f;
mem[2108] = 8'h3f;
mem[2109] = 8'h3f;
mem[2110] = 8'h3f;
mem[2111] = 8'h00;
mem[2112] = 8'h00;
mem[2113] = 8'hfc;
mem[2114] = 8'hfc;
mem[2115] = 8'hfc;
mem[2116] = 8'hfc;
mem[2117] = 8'hfc;
mem[2118] = 8'hfc;
mem[2119] = 8'h00;
mem[2120] = 8'h00;
mem[2121] = 8'h54;
mem[2122] = 8'h2a;
mem[2123] = 8'h54;
mem[2124] = 8'h2a;
mem[2125] = 8'h54;
mem[2126] = 8'h2a;
mem[2127] = 8'h00;
mem[2128] = 8'h00;
mem[2129] = 8'h00;
mem[2130] = 8'h18;
mem[2131] = 8'h3c;
mem[2132] = 8'h3c;
mem[2133] = 8'h7e;
mem[2134] = 8'h7e;
mem[2135] = 8'h7e;
mem[2136] = 8'h7e;
mem[2137] = 8'h7e;
mem[2138] = 8'h7e;
mem[2139] = 8'h3c;
mem[2140] = 8'h3c;
mem[2141] = 8'h18;
mem[2142] = 8'h00;
mem[2143] = 8'h00;
mem[2144] = 8'h07;
mem[2145] = 8'h1f;
mem[2146] = 8'h3f;
mem[2147] = 8'h7f;
mem[2148] = 8'h7f;
mem[2149] = 8'hff;
mem[2150] = 8'hff;
mem[2151] = 8'hff;
mem[2152] = 8'he0;
mem[2153] = 8'hf8;
mem[2154] = 8'hfc;
mem[2155] = 8'hfe;
mem[2156] = 8'hfe;
mem[2157] = 8'hff;
mem[2158] = 8'hff;
mem[2159] = 8'hff;
mem[2160] = 8'hff;
mem[2161] = 8'hff;
mem[2162] = 8'hff;
mem[2163] = 8'hfe;
mem[2164] = 8'hfe;
mem[2165] = 8'hfc;
mem[2166] = 8'hf8;
mem[2167] = 8'he0;
mem[2168] = 8'hff;
mem[2169] = 8'hff;
mem[2170] = 8'hff;
mem[2171] = 8'h7f;
mem[2172] = 8'h7f;
mem[2173] = 8'h3f;
mem[2174] = 8'h1f;
mem[2175] = 8'h07;
mem[2176] = 8'h24;
mem[2177] = 8'h42;
mem[2178] = 8'h81;
mem[2179] = 8'h00;
mem[2180] = 8'h00;
mem[2181] = 8'h81;
mem[2182] = 8'h42;
mem[2183] = 8'h24;
mem[2184] = 8'h00;
mem[2185] = 8'h00;
mem[2186] = 8'h02;
mem[2187] = 8'h00;
mem[2188] = 8'h00;
mem[2189] = 8'h00;
mem[2190] = 8'h20;
mem[2191] = 8'h00;
mem[2192] = 8'h20;
mem[2193] = 8'h00;
mem[2194] = 8'h02;
mem[2195] = 8'h00;
mem[2196] = 8'h20;
mem[2197] = 8'h00;
mem[2198] = 8'h02;
mem[2199] = 8'h00;
mem[2200] = 8'h22;
mem[2201] = 8'h00;
mem[2202] = 8'h88;
mem[2203] = 8'h00;
mem[2204] = 8'h22;
mem[2205] = 8'h00;
mem[2206] = 8'h88;
mem[2207] = 8'h00;
mem[2208] = 8'h88;
mem[2209] = 8'h00;
mem[2210] = 8'h55;
mem[2211] = 8'h00;
mem[2212] = 8'h22;
mem[2213] = 8'h00;
mem[2214] = 8'h55;
mem[2215] = 8'h00;
mem[2216] = 8'hff;
mem[2217] = 8'hbb;
mem[2218] = 8'hff;
mem[2219] = 8'hee;
mem[2220] = 8'hff;
mem[2221] = 8'hbb;
mem[2222] = 8'hff;
mem[2223] = 8'hee;
mem[2224] = 8'hbf;
mem[2225] = 8'hff;
mem[2226] = 8'hfb;
mem[2227] = 8'hff;
mem[2228] = 8'hbf;
mem[2229] = 8'hff;
mem[2230] = 8'hfb;
mem[2231] = 8'hff;
mem[2232] = 8'hff;
mem[2233] = 8'hff;
mem[2234] = 8'hdf;
mem[2235] = 8'hff;
mem[2236] = 8'hff;
mem[2237] = 8'hff;
mem[2238] = 8'hfd;
mem[2239] = 8'hff;
mem[2240] = 8'haa;
mem[2241] = 8'h00;
mem[2242] = 8'haa;
mem[2243] = 8'h00;
mem[2244] = 8'haa;
mem[2245] = 8'h00;
mem[2246] = 8'haa;
mem[2247] = 8'h00;
mem[2248] = 8'h00;
mem[2249] = 8'h44;
mem[2250] = 8'h00;
mem[2251] = 8'h00;
mem[2252] = 8'h00;
mem[2253] = 8'h44;
mem[2254] = 8'h00;
mem[2255] = 8'h00;
mem[2256] = 8'hcc;
mem[2257] = 8'hcc;
mem[2258] = 8'h33;
mem[2259] = 8'h33;
mem[2260] = 8'hcc;
mem[2261] = 8'hcc;
mem[2262] = 8'h33;
mem[2263] = 8'h33;
mem[2264] = 8'h3c;
mem[2265] = 8'h66;
mem[2266] = 8'h66;
mem[2267] = 8'h30;
mem[2268] = 8'h18;
mem[2269] = 8'h00;
mem[2270] = 8'h18;
mem[2271] = 8'h00;
mem[2272] = 8'h33;
mem[2273] = 8'h66;
mem[2274] = 8'hcc;
mem[2275] = 8'h99;
mem[2276] = 8'h33;
mem[2277] = 8'h66;
mem[2278] = 8'hcc;
mem[2279] = 8'h99;
mem[2280] = 8'hcc;
mem[2281] = 8'h66;
mem[2282] = 8'h33;
mem[2283] = 8'h99;
mem[2284] = 8'hcc;
mem[2285] = 8'h66;
mem[2286] = 8'h33;
mem[2287] = 8'h99;
mem[2288] = 8'he0;
mem[2289] = 8'ha0;
mem[2290] = 8'hee;
mem[2291] = 8'hc8;
mem[2292] = 8'hae;
mem[2293] = 8'h02;
mem[2294] = 8'h0e;
mem[2295] = 8'h00;
mem[2296] = 8'ha0;
mem[2297] = 8'ha0;
mem[2298] = 8'hae;
mem[2299] = 8'ha8;
mem[2300] = 8'hee;
mem[2301] = 8'h02;
mem[2302] = 8'h0e;
mem[2303] = 8'h00;
mem[2304] = 8'h00;
mem[2305] = 8'h00;
mem[2306] = 8'h00;
mem[2307] = 8'h00;
mem[2308] = 8'h00;
mem[2309] = 8'h00;
mem[2310] = 8'h00;
mem[2311] = 8'h00;
mem[2312] = 8'h18;
mem[2313] = 8'h18;
mem[2314] = 8'h18;
mem[2315] = 8'h18;
mem[2316] = 8'h18;
mem[2317] = 8'h00;
mem[2318] = 8'h18;
mem[2319] = 8'h00;
mem[2320] = 8'h66;
mem[2321] = 8'h66;
mem[2322] = 8'h66;
mem[2323] = 8'h00;
mem[2324] = 8'h00;
mem[2325] = 8'h00;
mem[2326] = 8'h00;
mem[2327] = 8'h00;
mem[2328] = 8'h6c;
mem[2329] = 8'h6c;
mem[2330] = 8'hfe;
mem[2331] = 8'h6c;
mem[2332] = 8'hfe;
mem[2333] = 8'h6c;
mem[2334] = 8'h6c;
mem[2335] = 8'h00;
mem[2336] = 8'h18;
mem[2337] = 8'h3e;
mem[2338] = 8'h60;
mem[2339] = 8'h3c;
mem[2340] = 8'h06;
mem[2341] = 8'h7c;
mem[2342] = 8'h18;
mem[2343] = 8'h00;
mem[2344] = 8'h00;
mem[2345] = 8'hc6;
mem[2346] = 8'hcc;
mem[2347] = 8'h18;
mem[2348] = 8'h30;
mem[2349] = 8'h66;
mem[2350] = 8'hc6;
mem[2351] = 8'h00;
mem[2352] = 8'h38;
mem[2353] = 8'h6c;
mem[2354] = 8'h38;
mem[2355] = 8'h76;
mem[2356] = 8'hdc;
mem[2357] = 8'hcc;
mem[2358] = 8'h76;
mem[2359] = 8'h00;
mem[2360] = 8'h18;
mem[2361] = 8'h18;
mem[2362] = 8'h30;
mem[2363] = 8'h00;
mem[2364] = 8'h00;
mem[2365] = 8'h00;
mem[2366] = 8'h00;
mem[2367] = 8'h00;
mem[2368] = 8'h0c;
mem[2369] = 8'h18;
mem[2370] = 8'h30;
mem[2371] = 8'h30;
mem[2372] = 8'h30;
mem[2373] = 8'h18;
mem[2374] = 8'h0c;
mem[2375] = 8'h00;
mem[2376] = 8'h30;
mem[2377] = 8'h18;
mem[2378] = 8'h0c;
mem[2379] = 8'h0c;
mem[2380] = 8'h0c;
mem[2381] = 8'h18;
mem[2382] = 8'h30;
mem[2383] = 8'h00;
mem[2384] = 8'h00;
mem[2385] = 8'h66;
mem[2386] = 8'h3c;
mem[2387] = 8'hff;
mem[2388] = 8'h3c;
mem[2389] = 8'h66;
mem[2390] = 8'h00;
mem[2391] = 8'h00;
mem[2392] = 8'h00;
mem[2393] = 8'h18;
mem[2394] = 8'h18;
mem[2395] = 8'h7e;
mem[2396] = 8'h18;
mem[2397] = 8'h18;
mem[2398] = 8'h00;
mem[2399] = 8'h00;
mem[2400] = 8'h00;
mem[2401] = 8'h00;
mem[2402] = 8'h00;
mem[2403] = 8'h00;
mem[2404] = 8'h00;
mem[2405] = 8'h18;
mem[2406] = 8'h18;
mem[2407] = 8'h30;
mem[2408] = 8'h00;
mem[2409] = 8'h00;
mem[2410] = 8'h00;
mem[2411] = 8'h7e;
mem[2412] = 8'h00;
mem[2413] = 8'h00;
mem[2414] = 8'h00;
mem[2415] = 8'h00;
mem[2416] = 8'h00;
mem[2417] = 8'h00;
mem[2418] = 8'h00;
mem[2419] = 8'h00;
mem[2420] = 8'h00;
mem[2421] = 8'h18;
mem[2422] = 8'h18;
mem[2423] = 8'h00;
mem[2424] = 8'h03;
mem[2425] = 8'h06;
mem[2426] = 8'h0c;
mem[2427] = 8'h18;
mem[2428] = 8'h30;
mem[2429] = 8'h60;
mem[2430] = 8'hc0;
mem[2431] = 8'h00;
mem[2432] = 8'h3c;
mem[2433] = 8'h66;
mem[2434] = 8'h6e;
mem[2435] = 8'h76;
mem[2436] = 8'h66;
mem[2437] = 8'h66;
mem[2438] = 8'h3c;
mem[2439] = 8'h00;
mem[2440] = 8'h18;
mem[2441] = 8'h38;
mem[2442] = 8'h18;
mem[2443] = 8'h18;
mem[2444] = 8'h18;
mem[2445] = 8'h18;
mem[2446] = 8'h7e;
mem[2447] = 8'h00;
mem[2448] = 8'h3c;
mem[2449] = 8'h66;
mem[2450] = 8'h0c;
mem[2451] = 8'h18;
mem[2452] = 8'h30;
mem[2453] = 8'h60;
mem[2454] = 8'h7e;
mem[2455] = 8'h00;
mem[2456] = 8'h3c;
mem[2457] = 8'h66;
mem[2458] = 8'h06;
mem[2459] = 8'h1c;
mem[2460] = 8'h06;
mem[2461] = 8'h66;
mem[2462] = 8'h3c;
mem[2463] = 8'h00;
mem[2464] = 8'h1c;
mem[2465] = 8'h3c;
mem[2466] = 8'h6c;
mem[2467] = 8'hcc;
mem[2468] = 8'hfe;
mem[2469] = 8'h0c;
mem[2470] = 8'h0c;
mem[2471] = 8'h00;
mem[2472] = 8'h7e;
mem[2473] = 8'h60;
mem[2474] = 8'h7c;
mem[2475] = 8'h06;
mem[2476] = 8'h06;
mem[2477] = 8'h66;
mem[2478] = 8'h3c;
mem[2479] = 8'h00;
mem[2480] = 8'h1c;
mem[2481] = 8'h30;
mem[2482] = 8'h60;
mem[2483] = 8'h7c;
mem[2484] = 8'h66;
mem[2485] = 8'h66;
mem[2486] = 8'h3c;
mem[2487] = 8'h00;
mem[2488] = 8'h7e;
mem[2489] = 8'h06;
mem[2490] = 8'h06;
mem[2491] = 8'h0c;
mem[2492] = 8'h18;
mem[2493] = 8'h18;
mem[2494] = 8'h18;
mem[2495] = 8'h00;
mem[2496] = 8'h3c;
mem[2497] = 8'h66;
mem[2498] = 8'h66;
mem[2499] = 8'h3c;
mem[2500] = 8'h66;
mem[2501] = 8'h66;
mem[2502] = 8'h3c;
mem[2503] = 8'h00;
mem[2504] = 8'h3c;
mem[2505] = 8'h66;
mem[2506] = 8'h66;
mem[2507] = 8'h3e;
mem[2508] = 8'h06;
mem[2509] = 8'h0c;
mem[2510] = 8'h38;
mem[2511] = 8'h00;
mem[2512] = 8'h00;
mem[2513] = 8'h18;
mem[2514] = 8'h18;
mem[2515] = 8'h00;
mem[2516] = 8'h00;
mem[2517] = 8'h18;
mem[2518] = 8'h18;
mem[2519] = 8'h00;
mem[2520] = 8'h00;
mem[2521] = 8'h18;
mem[2522] = 8'h18;
mem[2523] = 8'h00;
mem[2524] = 8'h00;
mem[2525] = 8'h18;
mem[2526] = 8'h18;
mem[2527] = 8'h30;
mem[2528] = 8'h0c;
mem[2529] = 8'h18;
mem[2530] = 8'h30;
mem[2531] = 8'h60;
mem[2532] = 8'h30;
mem[2533] = 8'h18;
mem[2534] = 8'h0c;
mem[2535] = 8'h00;
mem[2536] = 8'h00;
mem[2537] = 8'h00;
mem[2538] = 8'h7e;
mem[2539] = 8'h00;
mem[2540] = 8'h7e;
mem[2541] = 8'h00;
mem[2542] = 8'h00;
mem[2543] = 8'h00;
mem[2544] = 8'h60;
mem[2545] = 8'h30;
mem[2546] = 8'h18;
mem[2547] = 8'h0c;
mem[2548] = 8'h18;
mem[2549] = 8'h30;
mem[2550] = 8'h60;
mem[2551] = 8'h00;
mem[2552] = 8'h3c;
mem[2553] = 8'h66;
mem[2554] = 8'h06;
mem[2555] = 8'h0c;
mem[2556] = 8'h18;
mem[2557] = 8'h00;
mem[2558] = 8'h18;
mem[2559] = 8'h00;
mem[2560] = 8'h7c;
mem[2561] = 8'hc6;
mem[2562] = 8'hde;
mem[2563] = 8'hde;
mem[2564] = 8'hde;
mem[2565] = 8'hc0;
mem[2566] = 8'h7c;
mem[2567] = 8'h00;
mem[2568] = 8'h18;
mem[2569] = 8'h3c;
mem[2570] = 8'h66;
mem[2571] = 8'h66;
mem[2572] = 8'h7e;
mem[2573] = 8'h66;
mem[2574] = 8'h66;
mem[2575] = 8'h00;
mem[2576] = 8'h7c;
mem[2577] = 8'h66;
mem[2578] = 8'h66;
mem[2579] = 8'h7c;
mem[2580] = 8'h66;
mem[2581] = 8'h66;
mem[2582] = 8'h7c;
mem[2583] = 8'h00;
mem[2584] = 8'h3c;
mem[2585] = 8'h66;
mem[2586] = 8'h60;
mem[2587] = 8'h60;
mem[2588] = 8'h60;
mem[2589] = 8'h66;
mem[2590] = 8'h3c;
mem[2591] = 8'h00;
mem[2592] = 8'h78;
mem[2593] = 8'h6c;
mem[2594] = 8'h66;
mem[2595] = 8'h66;
mem[2596] = 8'h66;
mem[2597] = 8'h6c;
mem[2598] = 8'h78;
mem[2599] = 8'h00;
mem[2600] = 8'h7e;
mem[2601] = 8'h60;
mem[2602] = 8'h60;
mem[2603] = 8'h7c;
mem[2604] = 8'h60;
mem[2605] = 8'h60;
mem[2606] = 8'h7e;
mem[2607] = 8'h00;
mem[2608] = 8'h7e;
mem[2609] = 8'h60;
mem[2610] = 8'h60;
mem[2611] = 8'h7c;
mem[2612] = 8'h60;
mem[2613] = 8'h60;
mem[2614] = 8'h60;
mem[2615] = 8'h00;
mem[2616] = 8'h3c;
mem[2617] = 8'h66;
mem[2618] = 8'h60;
mem[2619] = 8'h6e;
mem[2620] = 8'h66;
mem[2621] = 8'h66;
mem[2622] = 8'h3e;
mem[2623] = 8'h00;
mem[2624] = 8'h66;
mem[2625] = 8'h66;
mem[2626] = 8'h66;
mem[2627] = 8'h7e;
mem[2628] = 8'h66;
mem[2629] = 8'h66;
mem[2630] = 8'h66;
mem[2631] = 8'h00;
mem[2632] = 8'h7e;
mem[2633] = 8'h18;
mem[2634] = 8'h18;
mem[2635] = 8'h18;
mem[2636] = 8'h18;
mem[2637] = 8'h18;
mem[2638] = 8'h7e;
mem[2639] = 8'h00;
mem[2640] = 8'h06;
mem[2641] = 8'h06;
mem[2642] = 8'h06;
mem[2643] = 8'h06;
mem[2644] = 8'h06;
mem[2645] = 8'h66;
mem[2646] = 8'h3c;
mem[2647] = 8'h00;
mem[2648] = 8'hc6;
mem[2649] = 8'hcc;
mem[2650] = 8'hd8;
mem[2651] = 8'hf0;
mem[2652] = 8'hd8;
mem[2653] = 8'hcc;
mem[2654] = 8'hc6;
mem[2655] = 8'h00;
mem[2656] = 8'h60;
mem[2657] = 8'h60;
mem[2658] = 8'h60;
mem[2659] = 8'h60;
mem[2660] = 8'h60;
mem[2661] = 8'h60;
mem[2662] = 8'h7e;
mem[2663] = 8'h00;
mem[2664] = 8'hc6;
mem[2665] = 8'hee;
mem[2666] = 8'hfe;
mem[2667] = 8'hd6;
mem[2668] = 8'hc6;
mem[2669] = 8'hc6;
mem[2670] = 8'hc6;
mem[2671] = 8'h00;
mem[2672] = 8'hc6;
mem[2673] = 8'he6;
mem[2674] = 8'hf6;
mem[2675] = 8'hde;
mem[2676] = 8'hce;
mem[2677] = 8'hc6;
mem[2678] = 8'hc6;
mem[2679] = 8'h00;
mem[2680] = 8'h3c;
mem[2681] = 8'h66;
mem[2682] = 8'h66;
mem[2683] = 8'h66;
mem[2684] = 8'h66;
mem[2685] = 8'h66;
mem[2686] = 8'h3c;
mem[2687] = 8'h00;
mem[2688] = 8'h7c;
mem[2689] = 8'h66;
mem[2690] = 8'h66;
mem[2691] = 8'h7c;
mem[2692] = 8'h60;
mem[2693] = 8'h60;
mem[2694] = 8'h60;
mem[2695] = 8'h00;
mem[2696] = 8'h3c;
mem[2697] = 8'h66;
mem[2698] = 8'h66;
mem[2699] = 8'h66;
mem[2700] = 8'h66;
mem[2701] = 8'h6c;
mem[2702] = 8'h36;
mem[2703] = 8'h00;
mem[2704] = 8'h7c;
mem[2705] = 8'h66;
mem[2706] = 8'h66;
mem[2707] = 8'h7c;
mem[2708] = 8'h6c;
mem[2709] = 8'h66;
mem[2710] = 8'h66;
mem[2711] = 8'h00;
mem[2712] = 8'h3c;
mem[2713] = 8'h66;
mem[2714] = 8'h60;
mem[2715] = 8'h3c;
mem[2716] = 8'h06;
mem[2717] = 8'h66;
mem[2718] = 8'h3c;
mem[2719] = 8'h00;
mem[2720] = 8'h7e;
mem[2721] = 8'h18;
mem[2722] = 8'h18;
mem[2723] = 8'h18;
mem[2724] = 8'h18;
mem[2725] = 8'h18;
mem[2726] = 8'h18;
mem[2727] = 8'h00;
mem[2728] = 8'h66;
mem[2729] = 8'h66;
mem[2730] = 8'h66;
mem[2731] = 8'h66;
mem[2732] = 8'h66;
mem[2733] = 8'h66;
mem[2734] = 8'h3c;
mem[2735] = 8'h00;
mem[2736] = 8'h66;
mem[2737] = 8'h66;
mem[2738] = 8'h66;
mem[2739] = 8'h66;
mem[2740] = 8'h66;
mem[2741] = 8'h3c;
mem[2742] = 8'h18;
mem[2743] = 8'h00;
mem[2744] = 8'hc6;
mem[2745] = 8'hc6;
mem[2746] = 8'hc6;
mem[2747] = 8'hd6;
mem[2748] = 8'hfe;
mem[2749] = 8'hee;
mem[2750] = 8'hc6;
mem[2751] = 8'h00;
mem[2752] = 8'hc3;
mem[2753] = 8'h66;
mem[2754] = 8'h3c;
mem[2755] = 8'h18;
mem[2756] = 8'h3c;
mem[2757] = 8'h66;
mem[2758] = 8'hc3;
mem[2759] = 8'h00;
mem[2760] = 8'hc3;
mem[2761] = 8'h66;
mem[2762] = 8'h3c;
mem[2763] = 8'h18;
mem[2764] = 8'h18;
mem[2765] = 8'h18;
mem[2766] = 8'h18;
mem[2767] = 8'h00;
mem[2768] = 8'h7e;
mem[2769] = 8'h06;
mem[2770] = 8'h0c;
mem[2771] = 8'h18;
mem[2772] = 8'h30;
mem[2773] = 8'h60;
mem[2774] = 8'h7e;
mem[2775] = 8'h00;
mem[2776] = 8'h3c;
mem[2777] = 8'h30;
mem[2778] = 8'h30;
mem[2779] = 8'h30;
mem[2780] = 8'h30;
mem[2781] = 8'h30;
mem[2782] = 8'h3c;
mem[2783] = 8'h00;
mem[2784] = 8'hc0;
mem[2785] = 8'h60;
mem[2786] = 8'h30;
mem[2787] = 8'h18;
mem[2788] = 8'h0c;
mem[2789] = 8'h06;
mem[2790] = 8'h03;
mem[2791] = 8'h00;
mem[2792] = 8'h3c;
mem[2793] = 8'h0c;
mem[2794] = 8'h0c;
mem[2795] = 8'h0c;
mem[2796] = 8'h0c;
mem[2797] = 8'h0c;
mem[2798] = 8'h3c;
mem[2799] = 8'h00;
mem[2800] = 8'h10;
mem[2801] = 8'h38;
mem[2802] = 8'h6c;
mem[2803] = 8'hc6;
mem[2804] = 8'h00;
mem[2805] = 8'h00;
mem[2806] = 8'h00;
mem[2807] = 8'h00;
mem[2808] = 8'h00;
mem[2809] = 8'h00;
mem[2810] = 8'h00;
mem[2811] = 8'h00;
mem[2812] = 8'h00;
mem[2813] = 8'h00;
mem[2814] = 8'h00;
mem[2815] = 8'hff;
mem[2816] = 8'h18;
mem[2817] = 8'h0c;
mem[2818] = 8'h06;
mem[2819] = 8'h00;
mem[2820] = 8'h00;
mem[2821] = 8'h00;
mem[2822] = 8'h00;
mem[2823] = 8'h00;
mem[2824] = 8'h00;
mem[2825] = 8'h00;
mem[2826] = 8'h3c;
mem[2827] = 8'h06;
mem[2828] = 8'h3e;
mem[2829] = 8'h66;
mem[2830] = 8'h3e;
mem[2831] = 8'h00;
mem[2832] = 8'h60;
mem[2833] = 8'h60;
mem[2834] = 8'h7c;
mem[2835] = 8'h66;
mem[2836] = 8'h66;
mem[2837] = 8'h66;
mem[2838] = 8'h7c;
mem[2839] = 8'h00;
mem[2840] = 8'h00;
mem[2841] = 8'h00;
mem[2842] = 8'h3c;
mem[2843] = 8'h60;
mem[2844] = 8'h60;
mem[2845] = 8'h60;
mem[2846] = 8'h3c;
mem[2847] = 8'h00;
mem[2848] = 8'h06;
mem[2849] = 8'h06;
mem[2850] = 8'h3e;
mem[2851] = 8'h66;
mem[2852] = 8'h66;
mem[2853] = 8'h66;
mem[2854] = 8'h3e;
mem[2855] = 8'h00;
mem[2856] = 8'h00;
mem[2857] = 8'h00;
mem[2858] = 8'h3c;
mem[2859] = 8'h66;
mem[2860] = 8'h7e;
mem[2861] = 8'h60;
mem[2862] = 8'h3c;
mem[2863] = 8'h00;
mem[2864] = 8'h1c;
mem[2865] = 8'h30;
mem[2866] = 8'h7c;
mem[2867] = 8'h30;
mem[2868] = 8'h30;
mem[2869] = 8'h30;
mem[2870] = 8'h30;
mem[2871] = 8'h00;
mem[2872] = 8'h00;
mem[2873] = 8'h00;
mem[2874] = 8'h3e;
mem[2875] = 8'h66;
mem[2876] = 8'h66;
mem[2877] = 8'h3e;
mem[2878] = 8'h06;
mem[2879] = 8'h7c;
mem[2880] = 8'h60;
mem[2881] = 8'h60;
mem[2882] = 8'h7c;
mem[2883] = 8'h66;
mem[2884] = 8'h66;
mem[2885] = 8'h66;
mem[2886] = 8'h66;
mem[2887] = 8'h00;
mem[2888] = 8'h18;
mem[2889] = 8'h00;
mem[2890] = 8'h38;
mem[2891] = 8'h18;
mem[2892] = 8'h18;
mem[2893] = 8'h18;
mem[2894] = 8'h1e;
mem[2895] = 8'h00;
mem[2896] = 8'h0c;
mem[2897] = 8'h00;
mem[2898] = 8'h0c;
mem[2899] = 8'h0c;
mem[2900] = 8'h0c;
mem[2901] = 8'h0c;
mem[2902] = 8'h0c;
mem[2903] = 8'h78;
mem[2904] = 8'h60;
mem[2905] = 8'h60;
mem[2906] = 8'h66;
mem[2907] = 8'h6c;
mem[2908] = 8'h78;
mem[2909] = 8'h6c;
mem[2910] = 8'h66;
mem[2911] = 8'h00;
mem[2912] = 8'h38;
mem[2913] = 8'h18;
mem[2914] = 8'h18;
mem[2915] = 8'h18;
mem[2916] = 8'h18;
mem[2917] = 8'h18;
mem[2918] = 8'h1e;
mem[2919] = 8'h00;
mem[2920] = 8'h00;
mem[2921] = 8'h00;
mem[2922] = 8'hcc;
mem[2923] = 8'hfe;
mem[2924] = 8'hd6;
mem[2925] = 8'hd6;
mem[2926] = 8'hc6;
mem[2927] = 8'h00;
mem[2928] = 8'h00;
mem[2929] = 8'h00;
mem[2930] = 8'h7c;
mem[2931] = 8'h66;
mem[2932] = 8'h66;
mem[2933] = 8'h66;
mem[2934] = 8'h66;
mem[2935] = 8'h00;
mem[2936] = 8'h00;
mem[2937] = 8'h00;
mem[2938] = 8'h3c;
mem[2939] = 8'h66;
mem[2940] = 8'h66;
mem[2941] = 8'h66;
mem[2942] = 8'h3c;
mem[2943] = 8'h00;
mem[2944] = 8'h00;
mem[2945] = 8'h00;
mem[2946] = 8'h7c;
mem[2947] = 8'h66;
mem[2948] = 8'h66;
mem[2949] = 8'h7c;
mem[2950] = 8'h60;
mem[2951] = 8'h60;
mem[2952] = 8'h00;
mem[2953] = 8'h00;
mem[2954] = 8'h3e;
mem[2955] = 8'h66;
mem[2956] = 8'h66;
mem[2957] = 8'h3e;
mem[2958] = 8'h06;
mem[2959] = 8'h06;
mem[2960] = 8'h00;
mem[2961] = 8'h00;
mem[2962] = 8'h7c;
mem[2963] = 8'h66;
mem[2964] = 8'h60;
mem[2965] = 8'h60;
mem[2966] = 8'h60;
mem[2967] = 8'h00;
mem[2968] = 8'h00;
mem[2969] = 8'h00;
mem[2970] = 8'h3e;
mem[2971] = 8'h60;
mem[2972] = 8'h3c;
mem[2973] = 8'h06;
mem[2974] = 8'h7c;
mem[2975] = 8'h00;
mem[2976] = 8'h30;
mem[2977] = 8'h30;
mem[2978] = 8'h7e;
mem[2979] = 8'h30;
mem[2980] = 8'h30;
mem[2981] = 8'h30;
mem[2982] = 8'h1e;
mem[2983] = 8'h00;
mem[2984] = 8'h00;
mem[2985] = 8'h00;
mem[2986] = 8'h66;
mem[2987] = 8'h66;
mem[2988] = 8'h66;
mem[2989] = 8'h66;
mem[2990] = 8'h3e;
mem[2991] = 8'h00;
mem[2992] = 8'h00;
mem[2993] = 8'h00;
mem[2994] = 8'h66;
mem[2995] = 8'h66;
mem[2996] = 8'h66;
mem[2997] = 8'h3c;
mem[2998] = 8'h18;
mem[2999] = 8'h00;
mem[3000] = 8'h00;
mem[3001] = 8'h00;
mem[3002] = 8'hc6;
mem[3003] = 8'hc6;
mem[3004] = 8'hd6;
mem[3005] = 8'h7c;
mem[3006] = 8'h6c;
mem[3007] = 8'h00;
mem[3008] = 8'h00;
mem[3009] = 8'h00;
mem[3010] = 8'hc6;
mem[3011] = 8'h6c;
mem[3012] = 8'h38;
mem[3013] = 8'h6c;
mem[3014] = 8'hc6;
mem[3015] = 8'h00;
mem[3016] = 8'h00;
mem[3017] = 8'h00;
mem[3018] = 8'h66;
mem[3019] = 8'h66;
mem[3020] = 8'h66;
mem[3021] = 8'h3e;
mem[3022] = 8'h06;
mem[3023] = 8'h3c;
mem[3024] = 8'h00;
mem[3025] = 8'h00;
mem[3026] = 8'h7e;
mem[3027] = 8'h0c;
mem[3028] = 8'h18;
mem[3029] = 8'h30;
mem[3030] = 8'h7e;
mem[3031] = 8'h00;
mem[3032] = 8'h0e;
mem[3033] = 8'h18;
mem[3034] = 8'h18;
mem[3035] = 8'h70;
mem[3036] = 8'h18;
mem[3037] = 8'h18;
mem[3038] = 8'h0e;
mem[3039] = 8'h00;
mem[3040] = 8'h18;
mem[3041] = 8'h18;
mem[3042] = 8'h18;
mem[3043] = 8'h18;
mem[3044] = 8'h18;
mem[3045] = 8'h18;
mem[3046] = 8'h18;
mem[3047] = 8'h00;
mem[3048] = 8'h70;
mem[3049] = 8'h18;
mem[3050] = 8'h18;
mem[3051] = 8'h0e;
mem[3052] = 8'h18;
mem[3053] = 8'h18;
mem[3054] = 8'h70;
mem[3055] = 8'h00;
mem[3056] = 8'h76;
mem[3057] = 8'hdc;
mem[3058] = 8'h00;
mem[3059] = 8'h00;
mem[3060] = 8'h00;
mem[3061] = 8'h00;
mem[3062] = 8'h00;
mem[3063] = 8'h00;
mem[3064] = 8'hc0;
mem[3065] = 8'ha0;
mem[3066] = 8'hae;
mem[3067] = 8'ha4;
mem[3068] = 8'hc4;
mem[3069] = 8'h04;
mem[3070] = 8'h04;
mem[3071] = 8'h00;
mem[3072] = 8'h03;
mem[3073] = 8'h03;
mem[3074] = 8'h03;
mem[3075] = 8'h03;
mem[3076] = 8'h03;
mem[3077] = 8'h03;
mem[3078] = 8'h03;
mem[3079] = 8'h03;
mem[3080] = 8'h07;
mem[3081] = 8'h07;
mem[3082] = 8'h07;
mem[3083] = 8'h07;
mem[3084] = 8'h07;
mem[3085] = 8'h07;
mem[3086] = 8'h07;
mem[3087] = 8'h07;
mem[3088] = 8'h1f;
mem[3089] = 8'h1f;
mem[3090] = 8'h1f;
mem[3091] = 8'h1f;
mem[3092] = 8'h1f;
mem[3093] = 8'h1f;
mem[3094] = 8'h1f;
mem[3095] = 8'h1f;
mem[3096] = 8'h3f;
mem[3097] = 8'h3f;
mem[3098] = 8'h3f;
mem[3099] = 8'h3f;
mem[3100] = 8'h3f;
mem[3101] = 8'h3f;
mem[3102] = 8'h3f;
mem[3103] = 8'h3f;
mem[3104] = 8'h7f;
mem[3105] = 8'h7f;
mem[3106] = 8'h7f;
mem[3107] = 8'h7f;
mem[3108] = 8'h7f;
mem[3109] = 8'h7f;
mem[3110] = 8'h7f;
mem[3111] = 8'h7f;
mem[3112] = 8'hff;
mem[3113] = 8'hff;
mem[3114] = 8'h00;
mem[3115] = 8'h00;
mem[3116] = 8'h00;
mem[3117] = 8'h00;
mem[3118] = 8'h00;
mem[3119] = 8'h00;
mem[3120] = 8'hff;
mem[3121] = 8'hff;
mem[3122] = 8'hff;
mem[3123] = 8'h00;
mem[3124] = 8'h00;
mem[3125] = 8'h00;
mem[3126] = 8'h00;
mem[3127] = 8'h00;
mem[3128] = 8'hff;
mem[3129] = 8'hff;
mem[3130] = 8'hff;
mem[3131] = 8'hff;
mem[3132] = 8'hff;
mem[3133] = 8'h00;
mem[3134] = 8'h00;
mem[3135] = 8'h00;
mem[3136] = 8'hff;
mem[3137] = 8'hff;
mem[3138] = 8'hff;
mem[3139] = 8'hff;
mem[3140] = 8'hff;
mem[3141] = 8'hff;
mem[3142] = 8'h00;
mem[3143] = 8'h00;
mem[3144] = 8'hff;
mem[3145] = 8'hff;
mem[3146] = 8'hff;
mem[3147] = 8'hff;
mem[3148] = 8'hff;
mem[3149] = 8'hff;
mem[3150] = 8'hff;
mem[3151] = 8'h00;
mem[3152] = 8'haa;
mem[3153] = 8'h55;
mem[3154] = 8'haa;
mem[3155] = 8'h55;
mem[3156] = 8'h00;
mem[3157] = 8'h00;
mem[3158] = 8'h00;
mem[3159] = 8'h00;
mem[3160] = 8'h00;
mem[3161] = 8'h00;
mem[3162] = 8'h00;
mem[3163] = 8'h00;
mem[3164] = 8'haa;
mem[3165] = 8'h55;
mem[3166] = 8'haa;
mem[3167] = 8'h55;
mem[3168] = 8'ha0;
mem[3169] = 8'h50;
mem[3170] = 8'ha0;
mem[3171] = 8'h50;
mem[3172] = 8'ha0;
mem[3173] = 8'h50;
mem[3174] = 8'ha0;
mem[3175] = 8'h50;
mem[3176] = 8'h0a;
mem[3177] = 8'h05;
mem[3178] = 8'h0a;
mem[3179] = 8'h05;
mem[3180] = 8'h0a;
mem[3181] = 8'h05;
mem[3182] = 8'h0a;
mem[3183] = 8'h05;
mem[3184] = 8'hcc;
mem[3185] = 8'hcc;
mem[3186] = 8'h33;
mem[3187] = 8'h33;
mem[3188] = 8'h00;
mem[3189] = 8'h00;
mem[3190] = 8'h00;
mem[3191] = 8'h00;
mem[3192] = 8'h00;
mem[3193] = 8'h00;
mem[3194] = 8'h00;
mem[3195] = 8'h00;
mem[3196] = 8'hcc;
mem[3197] = 8'hcc;
mem[3198] = 8'h33;
mem[3199] = 8'h33;
mem[3200] = 8'hc0;
mem[3201] = 8'hc0;
mem[3202] = 8'h30;
mem[3203] = 8'h30;
mem[3204] = 8'hc0;
mem[3205] = 8'hc0;
mem[3206] = 8'h30;
mem[3207] = 8'h30;
mem[3208] = 8'h0c;
mem[3209] = 8'h0c;
mem[3210] = 8'h03;
mem[3211] = 8'h03;
mem[3212] = 8'h0c;
mem[3213] = 8'h0c;
mem[3214] = 8'h03;
mem[3215] = 8'h03;
mem[3216] = 8'h00;
mem[3217] = 8'h01;
mem[3218] = 8'h02;
mem[3219] = 8'h05;
mem[3220] = 8'h0a;
mem[3221] = 8'h15;
mem[3222] = 8'h2a;
mem[3223] = 8'h55;
mem[3224] = 8'h00;
mem[3225] = 8'h80;
mem[3226] = 8'h40;
mem[3227] = 8'ha0;
mem[3228] = 8'h50;
mem[3229] = 8'ha8;
mem[3230] = 8'h54;
mem[3231] = 8'haa;
mem[3232] = 8'haa;
mem[3233] = 8'h54;
mem[3234] = 8'ha8;
mem[3235] = 8'h50;
mem[3236] = 8'ha0;
mem[3237] = 8'h40;
mem[3238] = 8'h80;
mem[3239] = 8'h00;
mem[3240] = 8'haa;
mem[3241] = 8'h55;
mem[3242] = 8'h2a;
mem[3243] = 8'h15;
mem[3244] = 8'h0a;
mem[3245] = 8'h05;
mem[3246] = 8'h02;
mem[3247] = 8'h01;
mem[3248] = 8'h00;
mem[3249] = 8'h00;
mem[3250] = 8'h01;
mem[3251] = 8'h03;
mem[3252] = 8'h0f;
mem[3253] = 8'h1f;
mem[3254] = 8'h3f;
mem[3255] = 8'h7f;
mem[3256] = 8'h00;
mem[3257] = 8'h00;
mem[3258] = 8'h80;
mem[3259] = 8'hc0;
mem[3260] = 8'hf0;
mem[3261] = 8'hf8;
mem[3262] = 8'hfc;
mem[3263] = 8'hfe;
mem[3264] = 8'hfe;
mem[3265] = 8'hfc;
mem[3266] = 8'hf8;
mem[3267] = 8'hf0;
mem[3268] = 8'hc0;
mem[3269] = 8'h80;
mem[3270] = 8'h00;
mem[3271] = 8'h00;
mem[3272] = 8'h7f;
mem[3273] = 8'h3f;
mem[3274] = 8'h1f;
mem[3275] = 8'h0f;
mem[3276] = 8'h03;
mem[3277] = 8'h01;
mem[3278] = 8'h00;
mem[3279] = 8'h00;
mem[3280] = 8'hff;
mem[3281] = 8'hff;
mem[3282] = 8'hfe;
mem[3283] = 8'hfc;
mem[3284] = 8'hf0;
mem[3285] = 8'he0;
mem[3286] = 8'hc0;
mem[3287] = 8'h80;
mem[3288] = 8'hff;
mem[3289] = 8'hff;
mem[3290] = 8'h7f;
mem[3291] = 8'h3f;
mem[3292] = 8'h0f;
mem[3293] = 8'h07;
mem[3294] = 8'h03;
mem[3295] = 8'h01;
mem[3296] = 8'h01;
mem[3297] = 8'h03;
mem[3298] = 8'h07;
mem[3299] = 8'h0f;
mem[3300] = 8'h3f;
mem[3301] = 8'h7f;
mem[3302] = 8'hff;
mem[3303] = 8'hff;
mem[3304] = 8'h80;
mem[3305] = 8'hc0;
mem[3306] = 8'he0;
mem[3307] = 8'hf0;
mem[3308] = 8'hfc;
mem[3309] = 8'hfe;
mem[3310] = 8'hff;
mem[3311] = 8'hff;
mem[3312] = 8'h00;
mem[3313] = 8'h00;
mem[3314] = 8'h00;
mem[3315] = 8'h00;
mem[3316] = 8'h03;
mem[3317] = 8'h0f;
mem[3318] = 8'h3f;
mem[3319] = 8'hff;
mem[3320] = 8'h00;
mem[3321] = 8'h00;
mem[3322] = 8'h00;
mem[3323] = 8'h00;
mem[3324] = 8'hc0;
mem[3325] = 8'hf0;
mem[3326] = 8'hfc;
mem[3327] = 8'hff;
mem[3328] = 8'hff;
mem[3329] = 8'hfc;
mem[3330] = 8'hf0;
mem[3331] = 8'hc0;
mem[3332] = 8'h00;
mem[3333] = 8'h00;
mem[3334] = 8'h00;
mem[3335] = 8'h00;
mem[3336] = 8'hff;
mem[3337] = 8'h3f;
mem[3338] = 8'h0f;
mem[3339] = 8'h03;
mem[3340] = 8'h00;
mem[3341] = 8'h00;
mem[3342] = 8'h00;
mem[3343] = 8'h00;
mem[3344] = 8'hff;
mem[3345] = 8'hff;
mem[3346] = 8'hff;
mem[3347] = 8'hff;
mem[3348] = 8'hfc;
mem[3349] = 8'hf0;
mem[3350] = 8'hc0;
mem[3351] = 8'h00;
mem[3352] = 8'hff;
mem[3353] = 8'hff;
mem[3354] = 8'hff;
mem[3355] = 8'hff;
mem[3356] = 8'h3f;
mem[3357] = 8'h0f;
mem[3358] = 8'h03;
mem[3359] = 8'h00;
mem[3360] = 8'h00;
mem[3361] = 8'h03;
mem[3362] = 8'h0f;
mem[3363] = 8'h3f;
mem[3364] = 8'hff;
mem[3365] = 8'hff;
mem[3366] = 8'hff;
mem[3367] = 8'hff;
mem[3368] = 8'h00;
mem[3369] = 8'hc0;
mem[3370] = 8'hf0;
mem[3371] = 8'hfc;
mem[3372] = 8'hff;
mem[3373] = 8'hff;
mem[3374] = 8'hff;
mem[3375] = 8'hff;
mem[3376] = 8'h01;
mem[3377] = 8'h01;
mem[3378] = 8'h03;
mem[3379] = 8'h03;
mem[3380] = 8'h07;
mem[3381] = 8'h07;
mem[3382] = 8'h0f;
mem[3383] = 8'h0f;
mem[3384] = 8'h80;
mem[3385] = 8'h80;
mem[3386] = 8'hc0;
mem[3387] = 8'hc0;
mem[3388] = 8'he0;
mem[3389] = 8'he0;
mem[3390] = 8'hf0;
mem[3391] = 8'hf0;
mem[3392] = 8'hf0;
mem[3393] = 8'hf0;
mem[3394] = 8'he0;
mem[3395] = 8'he0;
mem[3396] = 8'hc0;
mem[3397] = 8'hc0;
mem[3398] = 8'h80;
mem[3399] = 8'h80;
mem[3400] = 8'h0f;
mem[3401] = 8'h0f;
mem[3402] = 8'h07;
mem[3403] = 8'h07;
mem[3404] = 8'h03;
mem[3405] = 8'h03;
mem[3406] = 8'h01;
mem[3407] = 8'h01;
mem[3408] = 8'hfe;
mem[3409] = 8'hfe;
mem[3410] = 8'hfc;
mem[3411] = 8'hfc;
mem[3412] = 8'hf8;
mem[3413] = 8'hf8;
mem[3414] = 8'hf0;
mem[3415] = 8'hf0;
mem[3416] = 8'h7f;
mem[3417] = 8'h7f;
mem[3418] = 8'h3f;
mem[3419] = 8'h3f;
mem[3420] = 8'h1f;
mem[3421] = 8'h1f;
mem[3422] = 8'h0f;
mem[3423] = 8'h0f;
mem[3424] = 8'h0f;
mem[3425] = 8'h0f;
mem[3426] = 8'h1f;
mem[3427] = 8'h1f;
mem[3428] = 8'h3f;
mem[3429] = 8'h3f;
mem[3430] = 8'h7f;
mem[3431] = 8'h7f;
mem[3432] = 8'hf0;
mem[3433] = 8'hf0;
mem[3434] = 8'hf8;
mem[3435] = 8'hf8;
mem[3436] = 8'hfc;
mem[3437] = 8'hfc;
mem[3438] = 8'hfe;
mem[3439] = 8'hfe;
mem[3440] = 8'h00;
mem[3441] = 8'h00;
mem[3442] = 8'h00;
mem[3443] = 8'h00;
mem[3444] = 8'h00;
mem[3445] = 8'h03;
mem[3446] = 8'h1f;
mem[3447] = 8'hff;
mem[3448] = 8'h00;
mem[3449] = 8'h00;
mem[3450] = 8'h00;
mem[3451] = 8'h00;
mem[3452] = 8'h00;
mem[3453] = 8'hc0;
mem[3454] = 8'hf8;
mem[3455] = 8'hff;
mem[3456] = 8'hff;
mem[3457] = 8'hf8;
mem[3458] = 8'hc0;
mem[3459] = 8'h00;
mem[3460] = 8'h00;
mem[3461] = 8'h00;
mem[3462] = 8'h00;
mem[3463] = 8'h00;
mem[3464] = 8'hff;
mem[3465] = 8'h1f;
mem[3466] = 8'h03;
mem[3467] = 8'h00;
mem[3468] = 8'h00;
mem[3469] = 8'h00;
mem[3470] = 8'h00;
mem[3471] = 8'h00;
mem[3472] = 8'hff;
mem[3473] = 8'hff;
mem[3474] = 8'hff;
mem[3475] = 8'hff;
mem[3476] = 8'hff;
mem[3477] = 8'hfc;
mem[3478] = 8'he0;
mem[3479] = 8'h00;
mem[3480] = 8'hff;
mem[3481] = 8'hff;
mem[3482] = 8'hff;
mem[3483] = 8'hff;
mem[3484] = 8'hff;
mem[3485] = 8'h3f;
mem[3486] = 8'h07;
mem[3487] = 8'h00;
mem[3488] = 8'h00;
mem[3489] = 8'h07;
mem[3490] = 8'h3f;
mem[3491] = 8'hff;
mem[3492] = 8'hff;
mem[3493] = 8'hff;
mem[3494] = 8'hff;
mem[3495] = 8'hff;
mem[3496] = 8'h00;
mem[3497] = 8'he0;
mem[3498] = 8'hfc;
mem[3499] = 8'hff;
mem[3500] = 8'hff;
mem[3501] = 8'hff;
mem[3502] = 8'hff;
mem[3503] = 8'hff;
mem[3504] = 8'h00;
mem[3505] = 8'h00;
mem[3506] = 8'h01;
mem[3507] = 8'h03;
mem[3508] = 8'h03;
mem[3509] = 8'h07;
mem[3510] = 8'h0f;
mem[3511] = 8'h0f;
mem[3512] = 8'h00;
mem[3513] = 8'h00;
mem[3514] = 8'h80;
mem[3515] = 8'hc0;
mem[3516] = 8'hc0;
mem[3517] = 8'he0;
mem[3518] = 8'hf0;
mem[3519] = 8'hf0;
mem[3520] = 8'hf0;
mem[3521] = 8'hf0;
mem[3522] = 8'he0;
mem[3523] = 8'hc0;
mem[3524] = 8'hc0;
mem[3525] = 8'h80;
mem[3526] = 8'h00;
mem[3527] = 8'h00;
mem[3528] = 8'h0f;
mem[3529] = 8'h0f;
mem[3530] = 8'h07;
mem[3531] = 8'h03;
mem[3532] = 8'h03;
mem[3533] = 8'h01;
mem[3534] = 8'h00;
mem[3535] = 8'h00;
mem[3536] = 8'hff;
mem[3537] = 8'hff;
mem[3538] = 8'hfe;
mem[3539] = 8'hfc;
mem[3540] = 8'hfc;
mem[3541] = 8'hf8;
mem[3542] = 8'hf0;
mem[3543] = 8'hf0;
mem[3544] = 8'hff;
mem[3545] = 8'hff;
mem[3546] = 8'h7f;
mem[3547] = 8'h3f;
mem[3548] = 8'h3f;
mem[3549] = 8'h1f;
mem[3550] = 8'h0f;
mem[3551] = 8'h0f;
mem[3552] = 8'h0f;
mem[3553] = 8'h0f;
mem[3554] = 8'h1f;
mem[3555] = 8'h3f;
mem[3556] = 8'h3f;
mem[3557] = 8'h7f;
mem[3558] = 8'hff;
mem[3559] = 8'hff;
mem[3560] = 8'hf0;
mem[3561] = 8'hf0;
mem[3562] = 8'hf8;
mem[3563] = 8'hfc;
mem[3564] = 8'hfc;
mem[3565] = 8'hfe;
mem[3566] = 8'hff;
mem[3567] = 8'hff;
mem[3568] = 8'h00;
mem[3569] = 8'h00;
mem[3570] = 8'h00;
mem[3571] = 8'h00;
mem[3572] = 8'h01;
mem[3573] = 8'h03;
mem[3574] = 8'h07;
mem[3575] = 8'h0f;
mem[3576] = 8'h00;
mem[3577] = 8'h00;
mem[3578] = 8'h00;
mem[3579] = 8'h00;
mem[3580] = 8'h80;
mem[3581] = 8'hc0;
mem[3582] = 8'he0;
mem[3583] = 8'hf0;
mem[3584] = 8'hf0;
mem[3585] = 8'he0;
mem[3586] = 8'hc0;
mem[3587] = 8'h80;
mem[3588] = 8'h00;
mem[3589] = 8'h00;
mem[3590] = 8'h00;
mem[3591] = 8'h00;
mem[3592] = 8'h0f;
mem[3593] = 8'h07;
mem[3594] = 8'h03;
mem[3595] = 8'h01;
mem[3596] = 8'h00;
mem[3597] = 8'h00;
mem[3598] = 8'h00;
mem[3599] = 8'h00;
mem[3600] = 8'hff;
mem[3601] = 8'hff;
mem[3602] = 8'hff;
mem[3603] = 8'hff;
mem[3604] = 8'hfe;
mem[3605] = 8'hfc;
mem[3606] = 8'hf8;
mem[3607] = 8'hf0;
mem[3608] = 8'hff;
mem[3609] = 8'hff;
mem[3610] = 8'hff;
mem[3611] = 8'hff;
mem[3612] = 8'h7f;
mem[3613] = 8'h3f;
mem[3614] = 8'h1f;
mem[3615] = 8'h0f;
mem[3616] = 8'h0f;
mem[3617] = 8'h1f;
mem[3618] = 8'h3f;
mem[3619] = 8'h7f;
mem[3620] = 8'hff;
mem[3621] = 8'hff;
mem[3622] = 8'hff;
mem[3623] = 8'hff;
mem[3624] = 8'hf0;
mem[3625] = 8'hf8;
mem[3626] = 8'hfc;
mem[3627] = 8'hfe;
mem[3628] = 8'hff;
mem[3629] = 8'hff;
mem[3630] = 8'hff;
mem[3631] = 8'hff;
mem[3632] = 8'h00;
mem[3633] = 8'h00;
mem[3634] = 8'h00;
mem[3635] = 8'h00;
mem[3636] = 8'h03;
mem[3637] = 8'h07;
mem[3638] = 8'h0f;
mem[3639] = 8'h0f;
mem[3640] = 8'h00;
mem[3641] = 8'h00;
mem[3642] = 8'h00;
mem[3643] = 8'h00;
mem[3644] = 8'hc0;
mem[3645] = 8'he0;
mem[3646] = 8'hf0;
mem[3647] = 8'hf0;
mem[3648] = 8'hf0;
mem[3649] = 8'hf0;
mem[3650] = 8'he0;
mem[3651] = 8'hc0;
mem[3652] = 8'h00;
mem[3653] = 8'h00;
mem[3654] = 8'h00;
mem[3655] = 8'h00;
mem[3656] = 8'h0f;
mem[3657] = 8'h0f;
mem[3658] = 8'h07;
mem[3659] = 8'h03;
mem[3660] = 8'h00;
mem[3661] = 8'h00;
mem[3662] = 8'h00;
mem[3663] = 8'h00;
mem[3664] = 8'h00;
mem[3665] = 8'h00;
mem[3666] = 8'h00;
mem[3667] = 8'h00;
mem[3668] = 8'h00;
mem[3669] = 8'h01;
mem[3670] = 8'h03;
mem[3671] = 8'h07;
mem[3672] = 8'h00;
mem[3673] = 8'h00;
mem[3674] = 8'h00;
mem[3675] = 8'h00;
mem[3676] = 8'h00;
mem[3677] = 8'h80;
mem[3678] = 8'hc0;
mem[3679] = 8'he0;
mem[3680] = 8'he0;
mem[3681] = 8'hc0;
mem[3682] = 8'h80;
mem[3683] = 8'h00;
mem[3684] = 8'h00;
mem[3685] = 8'h00;
mem[3686] = 8'h00;
mem[3687] = 8'h00;
mem[3688] = 8'h07;
mem[3689] = 8'h03;
mem[3690] = 8'h01;
mem[3691] = 8'h00;
mem[3692] = 8'h00;
mem[3693] = 8'h00;
mem[3694] = 8'h00;
mem[3695] = 8'h00;
mem[3696] = 8'hff;
mem[3697] = 8'hff;
mem[3698] = 8'hff;
mem[3699] = 8'hff;
mem[3700] = 8'hff;
mem[3701] = 8'hfe;
mem[3702] = 8'hfc;
mem[3703] = 8'hf8;
mem[3704] = 8'hff;
mem[3705] = 8'hff;
mem[3706] = 8'hff;
mem[3707] = 8'hff;
mem[3708] = 8'hff;
mem[3709] = 8'h7f;
mem[3710] = 8'h3f;
mem[3711] = 8'h1f;
mem[3712] = 8'h1f;
mem[3713] = 8'h3f;
mem[3714] = 8'h7f;
mem[3715] = 8'hff;
mem[3716] = 8'hff;
mem[3717] = 8'hff;
mem[3718] = 8'hff;
mem[3719] = 8'hff;
mem[3720] = 8'hf8;
mem[3721] = 8'hfc;
mem[3722] = 8'hfe;
mem[3723] = 8'hff;
mem[3724] = 8'hff;
mem[3725] = 8'hff;
mem[3726] = 8'hff;
mem[3727] = 8'hff;
mem[3728] = 8'h00;
mem[3729] = 8'h00;
mem[3730] = 8'h00;
mem[3731] = 8'h03;
mem[3732] = 8'h3f;
mem[3733] = 8'hff;
mem[3734] = 8'hff;
mem[3735] = 8'hff;
mem[3736] = 8'h00;
mem[3737] = 8'h00;
mem[3738] = 8'h00;
mem[3739] = 8'hc0;
mem[3740] = 8'hfc;
mem[3741] = 8'hff;
mem[3742] = 8'hff;
mem[3743] = 8'hff;
mem[3744] = 8'hff;
mem[3745] = 8'hff;
mem[3746] = 8'hff;
mem[3747] = 8'hfc;
mem[3748] = 8'hc0;
mem[3749] = 8'h00;
mem[3750] = 8'h00;
mem[3751] = 8'h00;
mem[3752] = 8'hff;
mem[3753] = 8'hff;
mem[3754] = 8'hff;
mem[3755] = 8'h3f;
mem[3756] = 8'h03;
mem[3757] = 8'h00;
mem[3758] = 8'h00;
mem[3759] = 8'h00;
mem[3760] = 8'hef;
mem[3761] = 8'hef;
mem[3762] = 8'hc7;
mem[3763] = 8'hc7;
mem[3764] = 8'h83;
mem[3765] = 8'h83;
mem[3766] = 8'h01;
mem[3767] = 8'h01;
mem[3768] = 8'h3f;
mem[3769] = 8'h0f;
mem[3770] = 8'h03;
mem[3771] = 8'h00;
mem[3772] = 8'h03;
mem[3773] = 8'h0f;
mem[3774] = 8'h3f;
mem[3775] = 8'hff;
mem[3776] = 8'h01;
mem[3777] = 8'h01;
mem[3778] = 8'h83;
mem[3779] = 8'h83;
mem[3780] = 8'hc7;
mem[3781] = 8'hc7;
mem[3782] = 8'hef;
mem[3783] = 8'hef;
mem[3784] = 8'hfc;
mem[3785] = 8'hf0;
mem[3786] = 8'hc0;
mem[3787] = 8'h00;
mem[3788] = 8'hc0;
mem[3789] = 8'hf0;
mem[3790] = 8'hfc;
mem[3791] = 8'hff;
mem[3792] = 8'h00;
mem[3793] = 8'h00;
mem[3794] = 8'h00;
mem[3795] = 8'h00;
mem[3796] = 8'h10;
mem[3797] = 8'h38;
mem[3798] = 8'h7c;
mem[3799] = 8'hfe;
mem[3800] = 8'h80;
mem[3801] = 8'hc0;
mem[3802] = 8'he0;
mem[3803] = 8'hf0;
mem[3804] = 8'he0;
mem[3805] = 8'hc0;
mem[3806] = 8'h80;
mem[3807] = 8'h00;
mem[3808] = 8'hfe;
mem[3809] = 8'h7c;
mem[3810] = 8'h38;
mem[3811] = 8'h10;
mem[3812] = 8'h00;
mem[3813] = 8'h00;
mem[3814] = 8'h00;
mem[3815] = 8'h00;
mem[3816] = 8'h01;
mem[3817] = 8'h03;
mem[3818] = 8'h07;
mem[3819] = 8'h0f;
mem[3820] = 8'h07;
mem[3821] = 8'h03;
mem[3822] = 8'h01;
mem[3823] = 8'h00;
mem[3824] = 8'hff;
mem[3825] = 8'hff;
mem[3826] = 8'hff;
mem[3827] = 8'hff;
mem[3828] = 8'hef;
mem[3829] = 8'hc7;
mem[3830] = 8'h83;
mem[3831] = 8'h01;
mem[3832] = 8'h7f;
mem[3833] = 8'h3f;
mem[3834] = 8'h1f;
mem[3835] = 8'h0f;
mem[3836] = 8'h1f;
mem[3837] = 8'h3f;
mem[3838] = 8'h7f;
mem[3839] = 8'hff;
mem[3840] = 8'h01;
mem[3841] = 8'h83;
mem[3842] = 8'hc7;
mem[3843] = 8'hef;
mem[3844] = 8'hff;
mem[3845] = 8'hff;
mem[3846] = 8'hff;
mem[3847] = 8'hff;
mem[3848] = 8'hfe;
mem[3849] = 8'hfc;
mem[3850] = 8'hf8;
mem[3851] = 8'hf0;
mem[3852] = 8'hf8;
mem[3853] = 8'hfc;
mem[3854] = 8'hfe;
mem[3855] = 8'hff;
mem[3856] = 8'h18;
mem[3857] = 8'h3c;
mem[3858] = 8'h7e;
mem[3859] = 8'hff;
mem[3860] = 8'hff;
mem[3861] = 8'hff;
mem[3862] = 8'hff;
mem[3863] = 8'hff;
mem[3864] = 8'hf8;
mem[3865] = 8'hfc;
mem[3866] = 8'hfe;
mem[3867] = 8'hff;
mem[3868] = 8'hff;
mem[3869] = 8'hfe;
mem[3870] = 8'hfc;
mem[3871] = 8'hf8;
mem[3872] = 8'hff;
mem[3873] = 8'hff;
mem[3874] = 8'hff;
mem[3875] = 8'hff;
mem[3876] = 8'hff;
mem[3877] = 8'h7e;
mem[3878] = 8'h3c;
mem[3879] = 8'h18;
mem[3880] = 8'h1f;
mem[3881] = 8'h3f;
mem[3882] = 8'h7f;
mem[3883] = 8'hff;
mem[3884] = 8'hff;
mem[3885] = 8'h7f;
mem[3886] = 8'h3f;
mem[3887] = 8'h1f;
mem[3888] = 8'he7;
mem[3889] = 8'hc3;
mem[3890] = 8'h81;
mem[3891] = 8'h00;
mem[3892] = 8'h00;
mem[3893] = 8'h00;
mem[3894] = 8'h00;
mem[3895] = 8'h00;
mem[3896] = 8'h07;
mem[3897] = 8'h03;
mem[3898] = 8'h01;
mem[3899] = 8'h00;
mem[3900] = 8'h00;
mem[3901] = 8'h01;
mem[3902] = 8'h03;
mem[3903] = 8'h07;
mem[3904] = 8'h00;
mem[3905] = 8'h00;
mem[3906] = 8'h00;
mem[3907] = 8'h00;
mem[3908] = 8'h00;
mem[3909] = 8'h81;
mem[3910] = 8'hc3;
mem[3911] = 8'he7;
mem[3912] = 8'he0;
mem[3913] = 8'hc0;
mem[3914] = 8'h80;
mem[3915] = 8'h00;
mem[3916] = 8'h00;
mem[3917] = 8'h80;
mem[3918] = 8'hc0;
mem[3919] = 8'he0;
mem[3920] = 8'hff;
mem[3921] = 8'h7e;
mem[3922] = 8'h3c;
mem[3923] = 8'h18;
mem[3924] = 8'h18;
mem[3925] = 8'h3c;
mem[3926] = 8'h7e;
mem[3927] = 8'hff;
mem[3928] = 8'h81;
mem[3929] = 8'hc3;
mem[3930] = 8'he7;
mem[3931] = 8'hff;
mem[3932] = 8'hff;
mem[3933] = 8'he7;
mem[3934] = 8'hc3;
mem[3935] = 8'h81;
mem[3936] = 8'hff;
mem[3937] = 8'hff;
mem[3938] = 8'hc0;
mem[3939] = 8'hc0;
mem[3940] = 8'hc0;
mem[3941] = 8'hc0;
mem[3942] = 8'hc0;
mem[3943] = 8'hc0;
mem[3944] = 8'hff;
mem[3945] = 8'hff;
mem[3946] = 8'h03;
mem[3947] = 8'h03;
mem[3948] = 8'h03;
mem[3949] = 8'h03;
mem[3950] = 8'h03;
mem[3951] = 8'h03;
mem[3952] = 8'h03;
mem[3953] = 8'h03;
mem[3954] = 8'h03;
mem[3955] = 8'h03;
mem[3956] = 8'h03;
mem[3957] = 8'h03;
mem[3958] = 8'hff;
mem[3959] = 8'hff;
mem[3960] = 8'hc0;
mem[3961] = 8'hc0;
mem[3962] = 8'hc0;
mem[3963] = 8'hc0;
mem[3964] = 8'hc0;
mem[3965] = 8'hc0;
mem[3966] = 8'hff;
mem[3967] = 8'hff;
mem[3968] = 8'h00;
mem[3969] = 8'hff;
mem[3970] = 8'hff;
mem[3971] = 8'h00;
mem[3972] = 8'h00;
mem[3973] = 8'h00;
mem[3974] = 8'h00;
mem[3975] = 8'h00;
mem[3976] = 8'h00;
mem[3977] = 8'h00;
mem[3978] = 8'hff;
mem[3979] = 8'hff;
mem[3980] = 8'h00;
mem[3981] = 8'h00;
mem[3982] = 8'h00;
mem[3983] = 8'h00;
mem[3984] = 8'h00;
mem[3985] = 8'h00;
mem[3986] = 8'h00;
mem[3987] = 8'hff;
mem[3988] = 8'hff;
mem[3989] = 8'h00;
mem[3990] = 8'h00;
mem[3991] = 8'h00;
mem[3992] = 8'h00;
mem[3993] = 8'h00;
mem[3994] = 8'h00;
mem[3995] = 8'h00;
mem[3996] = 8'hff;
mem[3997] = 8'hff;
mem[3998] = 8'h00;
mem[3999] = 8'h00;
mem[4000] = 8'h00;
mem[4001] = 8'h00;
mem[4002] = 8'h00;
mem[4003] = 8'h00;
mem[4004] = 8'h00;
mem[4005] = 8'hff;
mem[4006] = 8'hff;
mem[4007] = 8'h00;
mem[4008] = 8'h60;
mem[4009] = 8'h60;
mem[4010] = 8'h60;
mem[4011] = 8'h60;
mem[4012] = 8'h60;
mem[4013] = 8'h60;
mem[4014] = 8'h60;
mem[4015] = 8'h60;
mem[4016] = 8'h30;
mem[4017] = 8'h30;
mem[4018] = 8'h30;
mem[4019] = 8'h30;
mem[4020] = 8'h30;
mem[4021] = 8'h30;
mem[4022] = 8'h30;
mem[4023] = 8'h30;
mem[4024] = 8'h0c;
mem[4025] = 8'h0c;
mem[4026] = 8'h0c;
mem[4027] = 8'h0c;
mem[4028] = 8'h0c;
mem[4029] = 8'h0c;
mem[4030] = 8'h0c;
mem[4031] = 8'h0c;
mem[4032] = 8'h06;
mem[4033] = 8'h06;
mem[4034] = 8'h06;
mem[4035] = 8'h06;
mem[4036] = 8'h06;
mem[4037] = 8'h06;
mem[4038] = 8'h06;
mem[4039] = 8'h06;
mem[4040] = 8'he0;
mem[4041] = 8'h38;
mem[4042] = 8'h0e;
mem[4043] = 8'h03;
mem[4044] = 8'h00;
mem[4045] = 8'h00;
mem[4046] = 8'h00;
mem[4047] = 8'h00;
mem[4048] = 8'h00;
mem[4049] = 8'h00;
mem[4050] = 8'h00;
mem[4051] = 8'h80;
mem[4052] = 8'he0;
mem[4053] = 8'h38;
mem[4054] = 8'h0e;
mem[4055] = 8'h03;
mem[4056] = 8'h00;
mem[4057] = 8'h00;
mem[4058] = 8'h00;
mem[4059] = 8'h01;
mem[4060] = 8'h07;
mem[4061] = 8'h1c;
mem[4062] = 8'h70;
mem[4063] = 8'hc0;
mem[4064] = 8'h07;
mem[4065] = 8'h1c;
mem[4066] = 8'h70;
mem[4067] = 8'hc0;
mem[4068] = 8'h00;
mem[4069] = 8'h00;
mem[4070] = 8'h00;
mem[4071] = 8'h00;
mem[4072] = 8'h80;
mem[4073] = 8'hc0;
mem[4074] = 8'hc0;
mem[4075] = 8'h60;
mem[4076] = 8'h60;
mem[4077] = 8'h30;
mem[4078] = 8'h30;
mem[4079] = 8'h18;
mem[4080] = 8'h18;
mem[4081] = 8'h0c;
mem[4082] = 8'h0c;
mem[4083] = 8'h06;
mem[4084] = 8'h06;
mem[4085] = 8'h03;
mem[4086] = 8'h03;
mem[4087] = 8'h01;
mem[4088] = 8'h18;
mem[4089] = 8'h30;
mem[4090] = 8'h30;
mem[4091] = 8'h60;
mem[4092] = 8'h60;
mem[4093] = 8'hc0;
mem[4094] = 8'hc0;
mem[4095] = 8'h80;
